.SUBCKT ActorSubckt NNIN1 NNIN2 NNIN3 NNIN4 NNIN5 NNIN6 NNIN7 NNIN8 NNIN9 NNIN10 NNIN11 NNIN12 NNIN13 NNIN14 NNIN15 NNIN16 NNIN17 NNIN18 NNIN19 NNOUT1

* LAYER 1: LINEAR
B1_1 L1_1 0 V=(V(NNIN1)*(-0.114165)+V(NNIN2)*(0.161748)+V(NNIN3)*(-0.193945)+V(NNIN4)*(0.201070)+V(NNIN5)*(0.070640)+V(NNIN6)*(2.059755)+V(NNIN7)*(1.090456)+V(NNIN8)*(1.276819)+V(NNIN9)*(0.626841)+V(NNIN10)*(0.642415)+V(NNIN11)*(0.073358)+V(NNIN12)*(-0.138243)+V(NNIN13)*(0.009260)+V(NNIN14)*(-0.007330)+V(NNIN15)*(-0.124777)+V(NNIN16)*(0.287745)+V(NNIN17)*(0.004955)+V(NNIN18)*(-0.110164)+V(NNIN19)*(0.058347)+(0.253910))
B1_2 L1_2 0 V=(V(NNIN1)*(0.106160)+V(NNIN2)*(0.154560)+V(NNIN3)*(-0.058837)+V(NNIN4)*(0.250518)+V(NNIN5)*(0.216628)+V(NNIN6)*(-1.674088)+V(NNIN7)*(-1.280336)+V(NNIN8)*(-1.175834)+V(NNIN9)*(-0.899666)+V(NNIN10)*(-0.867531)+V(NNIN11)*(0.142302)+V(NNIN12)*(0.119469)+V(NNIN13)*(0.125988)+V(NNIN14)*(0.105616)+V(NNIN15)*(-0.151881)+V(NNIN16)*(-0.148757)+V(NNIN17)*(0.381521)+V(NNIN18)*(0.303028)+V(NNIN19)*(-0.226211)+(0.208070))
B1_3 L1_3 0 V=(V(NNIN1)*(0.155568)+V(NNIN2)*(0.225487)+V(NNIN3)*(0.067225)+V(NNIN4)*(0.220303)+V(NNIN5)*(-0.003268)+V(NNIN6)*(1.530138)+V(NNIN7)*(0.885752)+V(NNIN8)*(0.962373)+V(NNIN9)*(0.465854)+V(NNIN10)*(0.611857)+V(NNIN11)*(0.236480)+V(NNIN12)*(0.271122)+V(NNIN13)*(0.432638)+V(NNIN14)*(0.186114)+V(NNIN15)*(0.360421)+V(NNIN16)*(0.076338)+V(NNIN17)*(-0.191961)+V(NNIN18)*(1.726694)+V(NNIN19)*(-0.089605)+(0.406359))
B1_4 L1_4 0 V=(V(NNIN1)*(0.065179)+V(NNIN2)*(0.305021)+V(NNIN3)*(0.048088)+V(NNIN4)*(0.246285)+V(NNIN5)*(0.044157)+V(NNIN6)*(-1.917416)+V(NNIN7)*(-1.444557)+V(NNIN8)*(-0.877293)+V(NNIN9)*(-0.657985)+V(NNIN10)*(-0.736570)+V(NNIN11)*(0.291707)+V(NNIN12)*(0.088448)+V(NNIN13)*(0.053435)+V(NNIN14)*(0.390162)+V(NNIN15)*(0.201510)+V(NNIN16)*(0.113558)+V(NNIN17)*(0.265973)+V(NNIN18)*(0.411459)+V(NNIN19)*(0.096870)+(0.155165))
B1_5 L1_5 0 V=(V(NNIN1)*(-0.028163)+V(NNIN2)*(0.149803)+V(NNIN3)*(-0.105346)+V(NNIN4)*(-0.035011)+V(NNIN5)*(-0.052522)+V(NNIN6)*(-1.047663)+V(NNIN7)*(-1.216216)+V(NNIN8)*(-1.362103)+V(NNIN9)*(-1.274414)+V(NNIN10)*(-1.166117)+V(NNIN11)*(-0.223455)+V(NNIN12)*(0.127963)+V(NNIN13)*(-0.083148)+V(NNIN14)*(0.070996)+V(NNIN15)*(0.147211)+V(NNIN16)*(0.301389)+V(NNIN17)*(0.166398)+V(NNIN18)*(-0.454368)+V(NNIN19)*(-0.012778)+(0.280780))
B1_6 L1_6 0 V=(V(NNIN1)*(0.201676)+V(NNIN2)*(0.096559)+V(NNIN3)*(-0.177280)+V(NNIN4)*(0.136017)+V(NNIN5)*(-0.058236)+V(NNIN6)*(-1.017563)+V(NNIN7)*(-0.942906)+V(NNIN8)*(-1.013858)+V(NNIN9)*(-0.908324)+V(NNIN10)*(-1.022393)+V(NNIN11)*(-0.044119)+V(NNIN12)*(-0.097866)+V(NNIN13)*(-0.063942)+V(NNIN14)*(-0.258553)+V(NNIN15)*(0.039485)+V(NNIN16)*(0.432263)+V(NNIN17)*(0.054633)+V(NNIN18)*(0.598301)+V(NNIN19)*(0.211151)+(0.147434))
B1_7 L1_7 0 V=(V(NNIN1)*(-0.008438)+V(NNIN2)*(0.052909)+V(NNIN3)*(0.022201)+V(NNIN4)*(0.060753)+V(NNIN5)*(-0.100531)+V(NNIN6)*(1.948704)+V(NNIN7)*(1.371158)+V(NNIN8)*(1.242682)+V(NNIN9)*(1.014841)+V(NNIN10)*(0.690017)+V(NNIN11)*(0.013172)+V(NNIN12)*(-0.121490)+V(NNIN13)*(0.070952)+V(NNIN14)*(-0.036764)+V(NNIN15)*(0.084944)+V(NNIN16)*(0.066850)+V(NNIN17)*(0.015851)+V(NNIN18)*(0.506564)+V(NNIN19)*(0.046335)+(0.249390))
B1_8 L1_8 0 V=(V(NNIN1)*(0.185542)+V(NNIN2)*(-0.101182)+V(NNIN3)*(0.287927)+V(NNIN4)*(0.200402)+V(NNIN5)*(0.219546)+V(NNIN6)*(-1.492036)+V(NNIN7)*(-1.009296)+V(NNIN8)*(-0.659153)+V(NNIN9)*(-0.560510)+V(NNIN10)*(-0.336476)+V(NNIN11)*(0.019539)+V(NNIN12)*(0.099498)+V(NNIN13)*(-0.020444)+V(NNIN14)*(-0.058755)+V(NNIN15)*(0.119281)+V(NNIN16)*(-0.006268)+V(NNIN17)*(-0.059586)+V(NNIN18)*(0.029218)+V(NNIN19)*(-0.186737)+(-0.022143))
B1_9 L1_9 0 V=(V(NNIN1)*(0.227583)+V(NNIN2)*(-0.068566)+V(NNIN3)*(0.226676)+V(NNIN4)*(0.006769)+V(NNIN5)*(-0.108666)+V(NNIN6)*(1.996603)+V(NNIN7)*(1.417610)+V(NNIN8)*(1.010934)+V(NNIN9)*(0.692548)+V(NNIN10)*(0.694986)+V(NNIN11)*(-0.154719)+V(NNIN12)*(0.166480)+V(NNIN13)*(0.112145)+V(NNIN14)*(-0.229875)+V(NNIN15)*(0.118705)+V(NNIN16)*(0.208914)+V(NNIN17)*(-0.095222)+V(NNIN18)*(0.159966)+V(NNIN19)*(0.037423)+(0.042389))
B1_10 L1_10 0 V=(V(NNIN1)*(0.280024)+V(NNIN2)*(-0.137973)+V(NNIN3)*(-0.019841)+V(NNIN4)*(0.140995)+V(NNIN5)*(0.127268)+V(NNIN6)*(-1.774235)+V(NNIN7)*(-1.036317)+V(NNIN8)*(-0.735848)+V(NNIN9)*(-0.469691)+V(NNIN10)*(-0.689591)+V(NNIN11)*(0.002233)+V(NNIN12)*(0.145836)+V(NNIN13)*(0.089704)+V(NNIN14)*(0.081291)+V(NNIN15)*(-0.071698)+V(NNIN16)*(0.056986)+V(NNIN17)*(0.001244)+V(NNIN18)*(-0.100177)+V(NNIN19)*(-0.133812)+(-0.034095))
B1_11 L1_11 0 V=(V(NNIN1)*(-0.131382)+V(NNIN2)*(-0.120516)+V(NNIN3)*(-0.189524)+V(NNIN4)*(0.201499)+V(NNIN5)*(0.221860)+V(NNIN6)*(-1.866005)+V(NNIN7)*(-1.428918)+V(NNIN8)*(-1.123147)+V(NNIN9)*(-0.957969)+V(NNIN10)*(-1.006796)+V(NNIN11)*(-0.049157)+V(NNIN12)*(-0.059529)+V(NNIN13)*(-0.171060)+V(NNIN14)*(0.034866)+V(NNIN15)*(0.087887)+V(NNIN16)*(0.352838)+V(NNIN17)*(0.210815)+V(NNIN18)*(-0.516776)+V(NNIN19)*(0.172191)+(0.080432))
B1_12 L1_12 0 V=(V(NNIN1)*(0.092218)+V(NNIN2)*(0.175729)+V(NNIN3)*(0.008230)+V(NNIN4)*(0.107847)+V(NNIN5)*(0.227278)+V(NNIN6)*(-1.859836)+V(NNIN7)*(-1.038642)+V(NNIN8)*(-0.930332)+V(NNIN9)*(-0.524285)+V(NNIN10)*(-0.424142)+V(NNIN11)*(0.329455)+V(NNIN12)*(0.107399)+V(NNIN13)*(0.269190)+V(NNIN14)*(0.322315)+V(NNIN15)*(0.351201)+V(NNIN16)*(0.206363)+V(NNIN17)*(0.185195)+V(NNIN18)*(-0.533978)+V(NNIN19)*(-0.088924)+(0.164881))
B1_13 L1_13 0 V=(V(NNIN1)*(-0.229673)+V(NNIN2)*(-0.160524)+V(NNIN3)*(-0.214567)+V(NNIN4)*(-0.014328)+V(NNIN5)*(-0.199332)+V(NNIN6)*(0.612319)+V(NNIN7)*(0.445635)+V(NNIN8)*(0.258539)+V(NNIN9)*(0.053950)+V(NNIN10)*(0.298466)+V(NNIN11)*(0.082465)+V(NNIN12)*(0.155860)+V(NNIN13)*(0.171223)+V(NNIN14)*(0.128103)+V(NNIN15)*(-0.027507)+V(NNIN16)*(0.329450)+V(NNIN17)*(-0.088522)+V(NNIN18)*(-3.747950)+V(NNIN19)*(-0.009344)+(-0.027862))
B1_14 L1_14 0 V=(V(NNIN1)*(-0.219537)+V(NNIN2)*(-0.076165)+V(NNIN3)*(0.017018)+V(NNIN4)*(-0.082570)+V(NNIN5)*(-0.251704)+V(NNIN6)*(1.875731)+V(NNIN7)*(1.076583)+V(NNIN8)*(0.859602)+V(NNIN9)*(0.805044)+V(NNIN10)*(0.620730)+V(NNIN11)*(-0.052536)+V(NNIN12)*(0.106108)+V(NNIN13)*(0.095052)+V(NNIN14)*(-0.140205)+V(NNIN15)*(-0.001431)+V(NNIN16)*(0.381084)+V(NNIN17)*(-0.232316)+V(NNIN18)*(0.544241)+V(NNIN19)*(-0.024154)+(0.165536))
B1_15 L1_15 0 V=(V(NNIN1)*(0.121503)+V(NNIN2)*(-0.212598)+V(NNIN3)*(-0.221119)+V(NNIN4)*(-0.088743)+V(NNIN5)*(-0.043956)+V(NNIN6)*(-2.234352)+V(NNIN7)*(-1.752074)+V(NNIN8)*(-1.745198)+V(NNIN9)*(-1.486982)+V(NNIN10)*(-1.367340)+V(NNIN11)*(0.108547)+V(NNIN12)*(0.107528)+V(NNIN13)*(0.067612)+V(NNIN14)*(0.032329)+V(NNIN15)*(0.084660)+V(NNIN16)*(0.255962)+V(NNIN17)*(0.039878)+V(NNIN18)*(0.025882)+V(NNIN19)*(0.043062)+(0.308802))
B1_16 L1_16 0 V=(V(NNIN1)*(0.208684)+V(NNIN2)*(0.204153)+V(NNIN3)*(0.216619)+V(NNIN4)*(0.019663)+V(NNIN5)*(-0.076687)+V(NNIN6)*(-1.085633)+V(NNIN7)*(-1.214084)+V(NNIN8)*(-0.750784)+V(NNIN9)*(-0.947411)+V(NNIN10)*(-1.084954)+V(NNIN11)*(0.095164)+V(NNIN12)*(-0.008123)+V(NNIN13)*(-0.029275)+V(NNIN14)*(0.210431)+V(NNIN15)*(0.165118)+V(NNIN16)*(0.380087)+V(NNIN17)*(0.179279)+V(NNIN18)*(2.389961)+V(NNIN19)*(-0.035974)+(0.108866))
B1_17 L1_17 0 V=(V(NNIN1)*(0.233961)+V(NNIN2)*(0.189529)+V(NNIN3)*(0.112089)+V(NNIN4)*(-0.096881)+V(NNIN5)*(-0.040611)+V(NNIN6)*(2.105502)+V(NNIN7)*(1.593700)+V(NNIN8)*(1.229177)+V(NNIN9)*(1.091754)+V(NNIN10)*(0.823907)+V(NNIN11)*(0.107804)+V(NNIN12)*(0.097088)+V(NNIN13)*(0.008330)+V(NNIN14)*(-0.175889)+V(NNIN15)*(0.099997)+V(NNIN16)*(0.327227)+V(NNIN17)*(-0.130135)+V(NNIN18)*(0.243226)+V(NNIN19)*(0.137389)+(0.314906))
B1_18 L1_18 0 V=(V(NNIN1)*(0.189762)+V(NNIN2)*(-0.134224)+V(NNIN3)*(0.166340)+V(NNIN4)*(0.073163)+V(NNIN5)*(0.106567)+V(NNIN6)*(2.089409)+V(NNIN7)*(1.133146)+V(NNIN8)*(1.245871)+V(NNIN9)*(0.640285)+V(NNIN10)*(0.605942)+V(NNIN11)*(-0.078302)+V(NNIN12)*(0.061609)+V(NNIN13)*(0.024606)+V(NNIN14)*(-0.097046)+V(NNIN15)*(0.158082)+V(NNIN16)*(0.322305)+V(NNIN17)*(-0.078659)+V(NNIN18)*(0.050294)+V(NNIN19)*(0.129283)+(0.298319))
B1_19 L1_19 0 V=(V(NNIN1)*(-0.059988)+V(NNIN2)*(0.185576)+V(NNIN3)*(0.070566)+V(NNIN4)*(0.173536)+V(NNIN5)*(0.065628)+V(NNIN6)*(0.161238)+V(NNIN7)*(0.273235)+V(NNIN8)*(0.420335)+V(NNIN9)*(0.476919)+V(NNIN10)*(0.557853)+V(NNIN11)*(0.064455)+V(NNIN12)*(-0.012175)+V(NNIN13)*(-0.174305)+V(NNIN14)*(-0.110207)+V(NNIN15)*(0.193199)+V(NNIN16)*(-0.229746)+V(NNIN17)*(0.017020)+V(NNIN18)*(-0.383044)+V(NNIN19)*(0.043501)+(-0.141010))
B1_20 L1_20 0 V=(V(NNIN1)*(-0.046954)+V(NNIN2)*(0.178236)+V(NNIN3)*(0.033016)+V(NNIN4)*(0.017466)+V(NNIN5)*(-0.010044)+V(NNIN6)*(2.168165)+V(NNIN7)*(1.694979)+V(NNIN8)*(1.266445)+V(NNIN9)*(1.226193)+V(NNIN10)*(0.863749)+V(NNIN11)*(0.151650)+V(NNIN12)*(-0.092891)+V(NNIN13)*(0.063872)+V(NNIN14)*(0.006646)+V(NNIN15)*(0.058459)+V(NNIN16)*(0.269223)+V(NNIN17)*(-0.166110)+V(NNIN18)*(-0.137257)+V(NNIN19)*(0.096071)+(0.290793))
B1_21 L1_21 0 V=(V(NNIN1)*(0.130126)+V(NNIN2)*(0.287617)+V(NNIN3)*(0.073652)+V(NNIN4)*(0.257714)+V(NNIN5)*(0.309869)+V(NNIN6)*(-1.787172)+V(NNIN7)*(-1.240866)+V(NNIN8)*(-0.964805)+V(NNIN9)*(-0.805731)+V(NNIN10)*(-0.802401)+V(NNIN11)*(0.140923)+V(NNIN12)*(0.159190)+V(NNIN13)*(0.173975)+V(NNIN14)*(-0.018667)+V(NNIN15)*(-0.178215)+V(NNIN16)*(-0.022070)+V(NNIN17)*(0.110990)+V(NNIN18)*(0.149349)+V(NNIN19)*(-0.175753)+(-0.088846))
B1_22 L1_22 0 V=(V(NNIN1)*(0.242636)+V(NNIN2)*(0.111363)+V(NNIN3)*(0.188449)+V(NNIN4)*(0.059527)+V(NNIN5)*(0.284318)+V(NNIN6)*(-1.744526)+V(NNIN7)*(-1.435969)+V(NNIN8)*(-0.871756)+V(NNIN9)*(-0.741844)+V(NNIN10)*(-0.758136)+V(NNIN11)*(0.303481)+V(NNIN12)*(0.205784)+V(NNIN13)*(0.362172)+V(NNIN14)*(0.224034)+V(NNIN15)*(0.265233)+V(NNIN16)*(0.045807)+V(NNIN17)*(0.192253)+V(NNIN18)*(0.290082)+V(NNIN19)*(0.058430)+(0.216745))
B1_23 L1_23 0 V=(V(NNIN1)*(0.062284)+V(NNIN2)*(0.002972)+V(NNIN3)*(0.086294)+V(NNIN4)*(-0.085245)+V(NNIN5)*(0.035434)+V(NNIN6)*(1.580656)+V(NNIN7)*(1.166181)+V(NNIN8)*(0.954246)+V(NNIN9)*(0.784485)+V(NNIN10)*(0.803167)+V(NNIN11)*(0.209082)+V(NNIN12)*(0.088558)+V(NNIN13)*(-0.064627)+V(NNIN14)*(-0.128596)+V(NNIN15)*(0.067585)+V(NNIN16)*(0.320100)+V(NNIN17)*(-0.158152)+V(NNIN18)*(0.142088)+V(NNIN19)*(-0.012347)+(0.279714))
B1_24 L1_24 0 V=(V(NNIN1)*(-0.166888)+V(NNIN2)*(-0.006530)+V(NNIN3)*(-0.138172)+V(NNIN4)*(0.072413)+V(NNIN5)*(0.100704)+V(NNIN6)*(0.221220)+V(NNIN7)*(-0.248994)+V(NNIN8)*(-0.212549)+V(NNIN9)*(-0.123608)+V(NNIN10)*(-0.300017)+V(NNIN11)*(0.030168)+V(NNIN12)*(0.026271)+V(NNIN13)*(0.296442)+V(NNIN14)*(0.221750)+V(NNIN15)*(0.213554)+V(NNIN16)*(0.196115)+V(NNIN17)*(0.064229)+V(NNIN18)*(0.264847)+V(NNIN19)*(0.097372)+(-0.004469))
B1_25 L1_25 0 V=(V(NNIN1)*(0.138354)+V(NNIN2)*(-0.195615)+V(NNIN3)*(-0.076998)+V(NNIN4)*(-0.200698)+V(NNIN5)*(0.188096)+V(NNIN6)*(-1.470528)+V(NNIN7)*(-1.172023)+V(NNIN8)*(-0.997365)+V(NNIN9)*(-1.140417)+V(NNIN10)*(-1.262862)+V(NNIN11)*(-0.117204)+V(NNIN12)*(0.173572)+V(NNIN13)*(-0.183302)+V(NNIN14)*(0.198197)+V(NNIN15)*(0.107754)+V(NNIN16)*(0.265984)+V(NNIN17)*(0.249489)+V(NNIN18)*(-0.065488)+V(NNIN19)*(0.072914)+(-0.044596))
B1_26 L1_26 0 V=(V(NNIN1)*(0.076203)+V(NNIN2)*(-0.070312)+V(NNIN3)*(0.063311)+V(NNIN4)*(0.260667)+V(NNIN5)*(-0.098406)+V(NNIN6)*(-1.952455)+V(NNIN7)*(-1.530133)+V(NNIN8)*(-1.026517)+V(NNIN9)*(-0.983931)+V(NNIN10)*(-1.003858)+V(NNIN11)*(0.081603)+V(NNIN12)*(0.166075)+V(NNIN13)*(0.211668)+V(NNIN14)*(0.036340)+V(NNIN15)*(0.198742)+V(NNIN16)*(0.331813)+V(NNIN17)*(0.368004)+V(NNIN18)*(1.348437)+V(NNIN19)*(0.133943)+(-0.086555))
B1_27 L1_27 0 V=(V(NNIN1)*(0.259590)+V(NNIN2)*(0.004773)+V(NNIN3)*(-0.080583)+V(NNIN4)*(0.022161)+V(NNIN5)*(-0.002757)+V(NNIN6)*(0.230455)+V(NNIN7)*(0.318918)+V(NNIN8)*(0.507779)+V(NNIN9)*(0.505138)+V(NNIN10)*(0.346142)+V(NNIN11)*(-0.049825)+V(NNIN12)*(0.052165)+V(NNIN13)*(-0.025183)+V(NNIN14)*(-0.073614)+V(NNIN15)*(0.144424)+V(NNIN16)*(-0.066305)+V(NNIN17)*(-0.223951)+V(NNIN18)*(-0.352501)+V(NNIN19)*(0.130967)+(-0.233768))
B1_28 L1_28 0 V=(V(NNIN1)*(0.373002)+V(NNIN2)*(0.251067)+V(NNIN3)*(0.320823)+V(NNIN4)*(0.038805)+V(NNIN5)*(0.345018)+V(NNIN6)*(-1.620281)+V(NNIN7)*(-0.907528)+V(NNIN8)*(-0.902579)+V(NNIN9)*(-0.424040)+V(NNIN10)*(-0.678404)+V(NNIN11)*(0.328249)+V(NNIN12)*(0.101437)+V(NNIN13)*(0.011315)+V(NNIN14)*(0.290475)+V(NNIN15)*(0.187543)+V(NNIN16)*(0.221622)+V(NNIN17)*(0.059658)+V(NNIN18)*(-0.167397)+V(NNIN19)*(-0.142580)+(0.162873))
B1_29 L1_29 0 V=(V(NNIN1)*(0.197359)+V(NNIN2)*(-0.079744)+V(NNIN3)*(-0.044160)+V(NNIN4)*(-0.140922)+V(NNIN5)*(-0.095751)+V(NNIN6)*(1.975538)+V(NNIN7)*(1.167377)+V(NNIN8)*(0.975684)+V(NNIN9)*(0.870341)+V(NNIN10)*(0.693914)+V(NNIN11)*(-0.003467)+V(NNIN12)*(0.081136)+V(NNIN13)*(-0.101301)+V(NNIN14)*(0.154392)+V(NNIN15)*(-0.169563)+V(NNIN16)*(0.380429)+V(NNIN17)*(-0.041656)+V(NNIN18)*(-0.306670)+V(NNIN19)*(0.039355)+(0.134825))
B1_30 L1_30 0 V=(V(NNIN1)*(0.041981)+V(NNIN2)*(0.184322)+V(NNIN3)*(-0.044187)+V(NNIN4)*(0.345801)+V(NNIN5)*(-0.061860)+V(NNIN6)*(1.535787)+V(NNIN7)*(1.314672)+V(NNIN8)*(0.868614)+V(NNIN9)*(0.598614)+V(NNIN10)*(0.534346)+V(NNIN11)*(0.001274)+V(NNIN12)*(-0.101208)+V(NNIN13)*(0.064918)+V(NNIN14)*(-0.081558)+V(NNIN15)*(0.091491)+V(NNIN16)*(0.259570)+V(NNIN17)*(-0.099452)+V(NNIN18)*(0.263572)+V(NNIN19)*(0.094603)+(0.248306))
B1_31 L1_31 0 V=(V(NNIN1)*(0.316330)+V(NNIN2)*(-0.121402)+V(NNIN3)*(-0.079757)+V(NNIN4)*(-0.137736)+V(NNIN5)*(0.098336)+V(NNIN6)*(1.425245)+V(NNIN7)*(1.193325)+V(NNIN8)*(0.598877)+V(NNIN9)*(0.767321)+V(NNIN10)*(0.376044)+V(NNIN11)*(0.627037)+V(NNIN12)*(0.230220)+V(NNIN13)*(0.356359)+V(NNIN14)*(0.143221)+V(NNIN15)*(0.132972)+V(NNIN16)*(0.083154)+V(NNIN17)*(-0.132944)+V(NNIN18)*(-2.283550)+V(NNIN19)*(-0.208674)+(0.086825))
B1_32 L1_32 0 V=(V(NNIN1)*(0.245964)+V(NNIN2)*(0.145688)+V(NNIN3)*(0.194635)+V(NNIN4)*(0.213213)+V(NNIN5)*(0.095736)+V(NNIN6)*(-1.998479)+V(NNIN7)*(-1.558448)+V(NNIN8)*(-1.275386)+V(NNIN9)*(-0.774461)+V(NNIN10)*(-0.811898)+V(NNIN11)*(0.260433)+V(NNIN12)*(0.026437)+V(NNIN13)*(0.158908)+V(NNIN14)*(0.291524)+V(NNIN15)*(-0.006138)+V(NNIN16)*(-0.161614)+V(NNIN17)*(0.430397)+V(NNIN18)*(-0.030702)+V(NNIN19)*(0.037332)+(0.045913))
* ACTIVATION LAYER 1: RELU
B_ACT1_1 L_ACT1_1 0 V=(IF(V(L1_1)>0,V(L1_1),0))
B_ACT1_2 L_ACT1_2 0 V=(IF(V(L1_2)>0,V(L1_2),0))
B_ACT1_3 L_ACT1_3 0 V=(IF(V(L1_3)>0,V(L1_3),0))
B_ACT1_4 L_ACT1_4 0 V=(IF(V(L1_4)>0,V(L1_4),0))
B_ACT1_5 L_ACT1_5 0 V=(IF(V(L1_5)>0,V(L1_5),0))
B_ACT1_6 L_ACT1_6 0 V=(IF(V(L1_6)>0,V(L1_6),0))
B_ACT1_7 L_ACT1_7 0 V=(IF(V(L1_7)>0,V(L1_7),0))
B_ACT1_8 L_ACT1_8 0 V=(IF(V(L1_8)>0,V(L1_8),0))
B_ACT1_9 L_ACT1_9 0 V=(IF(V(L1_9)>0,V(L1_9),0))
B_ACT1_10 L_ACT1_10 0 V=(IF(V(L1_10)>0,V(L1_10),0))
B_ACT1_11 L_ACT1_11 0 V=(IF(V(L1_11)>0,V(L1_11),0))
B_ACT1_12 L_ACT1_12 0 V=(IF(V(L1_12)>0,V(L1_12),0))
B_ACT1_13 L_ACT1_13 0 V=(IF(V(L1_13)>0,V(L1_13),0))
B_ACT1_14 L_ACT1_14 0 V=(IF(V(L1_14)>0,V(L1_14),0))
B_ACT1_15 L_ACT1_15 0 V=(IF(V(L1_15)>0,V(L1_15),0))
B_ACT1_16 L_ACT1_16 0 V=(IF(V(L1_16)>0,V(L1_16),0))
B_ACT1_17 L_ACT1_17 0 V=(IF(V(L1_17)>0,V(L1_17),0))
B_ACT1_18 L_ACT1_18 0 V=(IF(V(L1_18)>0,V(L1_18),0))
B_ACT1_19 L_ACT1_19 0 V=(IF(V(L1_19)>0,V(L1_19),0))
B_ACT1_20 L_ACT1_20 0 V=(IF(V(L1_20)>0,V(L1_20),0))
B_ACT1_21 L_ACT1_21 0 V=(IF(V(L1_21)>0,V(L1_21),0))
B_ACT1_22 L_ACT1_22 0 V=(IF(V(L1_22)>0,V(L1_22),0))
B_ACT1_23 L_ACT1_23 0 V=(IF(V(L1_23)>0,V(L1_23),0))
B_ACT1_24 L_ACT1_24 0 V=(IF(V(L1_24)>0,V(L1_24),0))
B_ACT1_25 L_ACT1_25 0 V=(IF(V(L1_25)>0,V(L1_25),0))
B_ACT1_26 L_ACT1_26 0 V=(IF(V(L1_26)>0,V(L1_26),0))
B_ACT1_27 L_ACT1_27 0 V=(IF(V(L1_27)>0,V(L1_27),0))
B_ACT1_28 L_ACT1_28 0 V=(IF(V(L1_28)>0,V(L1_28),0))
B_ACT1_29 L_ACT1_29 0 V=(IF(V(L1_29)>0,V(L1_29),0))
B_ACT1_30 L_ACT1_30 0 V=(IF(V(L1_30)>0,V(L1_30),0))
B_ACT1_31 L_ACT1_31 0 V=(IF(V(L1_31)>0,V(L1_31),0))
B_ACT1_32 L_ACT1_32 0 V=(IF(V(L1_32)>0,V(L1_32),0))
* LAYER 2: LINEAR
B2_1 L2_1 0 V=(V(L_ACT1_1)*(0.020810)+V(L_ACT1_2)*(0.173981)+V(L_ACT1_3)*(-0.037384)+V(L_ACT1_4)*(0.088305)+V(L_ACT1_5)*(0.280282)+V(L_ACT1_6)*(0.259442)+V(L_ACT1_7)*(-0.217917)+V(L_ACT1_8)*(0.047484)+V(L_ACT1_9)*(0.137104)+V(L_ACT1_10)*(0.221393)+V(L_ACT1_11)*(0.190468)+V(L_ACT1_12)*(0.068395)+V(L_ACT1_13)*(-0.019815)+V(L_ACT1_14)*(-0.463553)+V(L_ACT1_15)*(0.239120)+V(L_ACT1_16)*(0.167244)+V(L_ACT1_17)*(0.114417)+V(L_ACT1_18)*(-0.121226)+V(L_ACT1_19)*(-0.040037)+V(L_ACT1_20)*(-0.049026)+V(L_ACT1_21)*(0.285778)+V(L_ACT1_22)*(0.220973)+V(L_ACT1_23)*(-0.097595)+V(L_ACT1_24)*(-0.195209)+V(L_ACT1_25)*(0.072457)+V(L_ACT1_26)*(0.259739)+V(L_ACT1_27)*(-0.089615)+V(L_ACT1_28)*(0.272208)+V(L_ACT1_29)*(-0.320898)+V(L_ACT1_30)*(0.043506)+V(L_ACT1_31)*(-0.033063)+V(L_ACT1_32)*(0.021228)+(0.053924))
B2_2 L2_2 0 V=(V(L_ACT1_1)*(-0.124028)+V(L_ACT1_2)*(0.304012)+V(L_ACT1_3)*(-0.219834)+V(L_ACT1_4)*(0.031305)+V(L_ACT1_5)*(0.237195)+V(L_ACT1_6)*(0.290460)+V(L_ACT1_7)*(-0.045422)+V(L_ACT1_8)*(0.085893)+V(L_ACT1_9)*(0.076160)+V(L_ACT1_10)*(0.148510)+V(L_ACT1_11)*(0.370183)+V(L_ACT1_12)*(0.329442)+V(L_ACT1_13)*(0.118235)+V(L_ACT1_14)*(-0.356061)+V(L_ACT1_15)*(0.379593)+V(L_ACT1_16)*(0.271443)+V(L_ACT1_17)*(0.136560)+V(L_ACT1_18)*(-0.035831)+V(L_ACT1_19)*(-0.205137)+V(L_ACT1_20)*(-0.031926)+V(L_ACT1_21)*(0.098084)+V(L_ACT1_22)*(0.029228)+V(L_ACT1_23)*(-0.017278)+V(L_ACT1_24)*(-0.078898)+V(L_ACT1_25)*(0.092770)+V(L_ACT1_26)*(0.114401)+V(L_ACT1_27)*(-0.193899)+V(L_ACT1_28)*(0.273323)+V(L_ACT1_29)*(-0.348800)+V(L_ACT1_30)*(-0.211344)+V(L_ACT1_31)*(-0.155361)+V(L_ACT1_32)*(0.319418)+(0.033128))
B2_3 L2_3 0 V=(V(L_ACT1_1)*(0.220176)+V(L_ACT1_2)*(-0.146424)+V(L_ACT1_3)*(-0.022592)+V(L_ACT1_4)*(-0.170171)+V(L_ACT1_5)*(0.025141)+V(L_ACT1_6)*(-0.051186)+V(L_ACT1_7)*(0.022040)+V(L_ACT1_8)*(0.088491)+V(L_ACT1_9)*(-0.065482)+V(L_ACT1_10)*(0.023890)+V(L_ACT1_11)*(-0.076379)+V(L_ACT1_12)*(0.104522)+V(L_ACT1_13)*(-0.000374)+V(L_ACT1_14)*(0.230070)+V(L_ACT1_15)*(-0.293275)+V(L_ACT1_16)*(-0.309838)+V(L_ACT1_17)*(-0.142026)+V(L_ACT1_18)*(0.174067)+V(L_ACT1_19)*(0.145664)+V(L_ACT1_20)*(-0.193976)+V(L_ACT1_21)*(0.115344)+V(L_ACT1_22)*(-0.134402)+V(L_ACT1_23)*(-0.019329)+V(L_ACT1_24)*(0.005805)+V(L_ACT1_25)*(0.023168)+V(L_ACT1_26)*(-0.435266)+V(L_ACT1_27)*(0.006174)+V(L_ACT1_28)*(-0.078257)+V(L_ACT1_29)*(0.041673)+V(L_ACT1_30)*(0.024907)+V(L_ACT1_31)*(0.219430)+V(L_ACT1_32)*(-0.111911)+(-0.157541))
B2_4 L2_4 0 V=(V(L_ACT1_1)*(0.186869)+V(L_ACT1_2)*(-0.062033)+V(L_ACT1_3)*(0.182494)+V(L_ACT1_4)*(0.179831)+V(L_ACT1_5)*(-0.062667)+V(L_ACT1_6)*(-0.104512)+V(L_ACT1_7)*(0.167369)+V(L_ACT1_8)*(-0.158455)+V(L_ACT1_9)*(0.152624)+V(L_ACT1_10)*(-0.017370)+V(L_ACT1_11)*(-0.083422)+V(L_ACT1_12)*(0.051418)+V(L_ACT1_13)*(-0.199409)+V(L_ACT1_14)*(0.465461)+V(L_ACT1_15)*(-0.077907)+V(L_ACT1_16)*(-0.041273)+V(L_ACT1_17)*(0.156210)+V(L_ACT1_18)*(0.149517)+V(L_ACT1_19)*(0.249050)+V(L_ACT1_20)*(0.302048)+V(L_ACT1_21)*(-0.234906)+V(L_ACT1_22)*(-0.063900)+V(L_ACT1_23)*(0.226074)+V(L_ACT1_24)*(-0.002225)+V(L_ACT1_25)*(-0.360078)+V(L_ACT1_26)*(0.058802)+V(L_ACT1_27)*(-0.103258)+V(L_ACT1_28)*(0.105469)+V(L_ACT1_29)*(0.304449)+V(L_ACT1_30)*(0.229281)+V(L_ACT1_31)*(0.031347)+V(L_ACT1_32)*(-0.138390)+(0.112670))
B2_5 L2_5 0 V=(V(L_ACT1_1)*(-0.123831)+V(L_ACT1_2)*(0.122656)+V(L_ACT1_3)*(0.338512)+V(L_ACT1_4)*(-0.133963)+V(L_ACT1_5)*(-0.274605)+V(L_ACT1_6)*(0.032534)+V(L_ACT1_7)*(0.177853)+V(L_ACT1_8)*(-0.046638)+V(L_ACT1_9)*(-0.108839)+V(L_ACT1_10)*(0.214735)+V(L_ACT1_11)*(-0.203280)+V(L_ACT1_12)*(0.069503)+V(L_ACT1_13)*(-0.061563)+V(L_ACT1_14)*(0.167091)+V(L_ACT1_15)*(-0.070282)+V(L_ACT1_16)*(0.014277)+V(L_ACT1_17)*(0.192649)+V(L_ACT1_18)*(0.013171)+V(L_ACT1_19)*(0.178290)+V(L_ACT1_20)*(0.054554)+V(L_ACT1_21)*(-0.100151)+V(L_ACT1_22)*(0.156627)+V(L_ACT1_23)*(0.086318)+V(L_ACT1_24)*(0.093037)+V(L_ACT1_25)*(-0.363544)+V(L_ACT1_26)*(0.097085)+V(L_ACT1_27)*(0.187539)+V(L_ACT1_28)*(0.174304)+V(L_ACT1_29)*(0.134694)+V(L_ACT1_30)*(-0.126019)+V(L_ACT1_31)*(0.292957)+V(L_ACT1_32)*(0.132905)+(-0.138439))
B2_6 L2_6 0 V=(V(L_ACT1_1)*(0.353470)+V(L_ACT1_2)*(-0.019530)+V(L_ACT1_3)*(0.316199)+V(L_ACT1_4)*(-0.124913)+V(L_ACT1_5)*(0.023068)+V(L_ACT1_6)*(0.095962)+V(L_ACT1_7)*(0.151473)+V(L_ACT1_8)*(-0.126917)+V(L_ACT1_9)*(0.252790)+V(L_ACT1_10)*(-0.022019)+V(L_ACT1_11)*(-0.249817)+V(L_ACT1_12)*(0.025245)+V(L_ACT1_13)*(-0.184228)+V(L_ACT1_14)*(0.578601)+V(L_ACT1_15)*(-0.165720)+V(L_ACT1_16)*(0.010343)+V(L_ACT1_17)*(0.356842)+V(L_ACT1_18)*(0.197257)+V(L_ACT1_19)*(0.129158)+V(L_ACT1_20)*(-0.014149)+V(L_ACT1_21)*(-0.115148)+V(L_ACT1_22)*(-0.000640)+V(L_ACT1_23)*(0.181629)+V(L_ACT1_24)*(-0.039287)+V(L_ACT1_25)*(-0.107158)+V(L_ACT1_26)*(-0.138941)+V(L_ACT1_27)*(0.145985)+V(L_ACT1_28)*(-0.127041)+V(L_ACT1_29)*(0.262127)+V(L_ACT1_30)*(0.185642)+V(L_ACT1_31)*(-0.023469)+V(L_ACT1_32)*(0.010389)+(0.151875))
B2_7 L2_7 0 V=(V(L_ACT1_1)*(0.099683)+V(L_ACT1_2)*(-0.135899)+V(L_ACT1_3)*(-0.075481)+V(L_ACT1_4)*(-0.081849)+V(L_ACT1_5)*(0.089708)+V(L_ACT1_6)*(0.037446)+V(L_ACT1_7)*(-0.129304)+V(L_ACT1_8)*(0.040971)+V(L_ACT1_9)*(-0.030334)+V(L_ACT1_10)*(0.100139)+V(L_ACT1_11)*(0.015607)+V(L_ACT1_12)*(-0.164285)+V(L_ACT1_13)*(-0.073297)+V(L_ACT1_14)*(0.029120)+V(L_ACT1_15)*(0.014010)+V(L_ACT1_16)*(-0.020938)+V(L_ACT1_17)*(0.082770)+V(L_ACT1_18)*(-0.072880)+V(L_ACT1_19)*(-0.020377)+V(L_ACT1_20)*(0.004940)+V(L_ACT1_21)*(-0.171527)+V(L_ACT1_22)*(-0.204212)+V(L_ACT1_23)*(0.123236)+V(L_ACT1_24)*(0.022144)+V(L_ACT1_25)*(-0.095107)+V(L_ACT1_26)*(0.124137)+V(L_ACT1_27)*(-0.159099)+V(L_ACT1_28)*(-0.023133)+V(L_ACT1_29)*(0.045073)+V(L_ACT1_30)*(-0.003210)+V(L_ACT1_31)*(0.116906)+V(L_ACT1_32)*(0.082684)+(-0.106810))
B2_8 L2_8 0 V=(V(L_ACT1_1)*(0.318581)+V(L_ACT1_2)*(-0.153041)+V(L_ACT1_3)*(0.313941)+V(L_ACT1_4)*(0.081804)+V(L_ACT1_5)*(0.097334)+V(L_ACT1_6)*(0.027762)+V(L_ACT1_7)*(0.417114)+V(L_ACT1_8)*(0.009279)+V(L_ACT1_9)*(0.165996)+V(L_ACT1_10)*(-0.104892)+V(L_ACT1_11)*(-0.194010)+V(L_ACT1_12)*(-0.061781)+V(L_ACT1_13)*(0.073456)+V(L_ACT1_14)*(0.418269)+V(L_ACT1_15)*(0.007042)+V(L_ACT1_16)*(0.177999)+V(L_ACT1_17)*(0.245011)+V(L_ACT1_18)*(0.269437)+V(L_ACT1_19)*(0.099431)+V(L_ACT1_20)*(0.103760)+V(L_ACT1_21)*(-0.072231)+V(L_ACT1_22)*(-0.086209)+V(L_ACT1_23)*(0.176900)+V(L_ACT1_24)*(0.070992)+V(L_ACT1_25)*(-0.215297)+V(L_ACT1_26)*(-0.154474)+V(L_ACT1_27)*(0.019845)+V(L_ACT1_28)*(-0.018974)+V(L_ACT1_29)*(0.493626)+V(L_ACT1_30)*(0.263640)+V(L_ACT1_31)*(0.073467)+V(L_ACT1_32)*(-0.225370)+(0.068193))
B2_9 L2_9 0 V=(V(L_ACT1_1)*(0.148932)+V(L_ACT1_2)*(-0.189292)+V(L_ACT1_3)*(0.252967)+V(L_ACT1_4)*(-0.177038)+V(L_ACT1_5)*(0.197758)+V(L_ACT1_6)*(-0.144249)+V(L_ACT1_7)*(0.112326)+V(L_ACT1_8)*(-0.160745)+V(L_ACT1_9)*(0.029598)+V(L_ACT1_10)*(-0.006093)+V(L_ACT1_11)*(0.019748)+V(L_ACT1_12)*(0.182854)+V(L_ACT1_13)*(0.650198)+V(L_ACT1_14)*(0.570649)+V(L_ACT1_15)*(0.385248)+V(L_ACT1_16)*(0.049743)+V(L_ACT1_17)*(0.240052)+V(L_ACT1_18)*(0.310348)+V(L_ACT1_19)*(-0.146855)+V(L_ACT1_20)*(0.221426)+V(L_ACT1_21)*(-0.341030)+V(L_ACT1_22)*(-0.170921)+V(L_ACT1_23)*(0.256935)+V(L_ACT1_24)*(0.266598)+V(L_ACT1_25)*(-0.384344)+V(L_ACT1_26)*(-0.243714)+V(L_ACT1_27)*(-0.155099)+V(L_ACT1_28)*(0.192506)+V(L_ACT1_29)*(0.320598)+V(L_ACT1_30)*(-0.042744)+V(L_ACT1_31)*(0.230090)+V(L_ACT1_32)*(-0.080504)+(0.040231))
B2_10 L2_10 0 V=(V(L_ACT1_1)*(0.038652)+V(L_ACT1_2)*(0.103105)+V(L_ACT1_3)*(0.313085)+V(L_ACT1_4)*(-0.025102)+V(L_ACT1_5)*(0.009149)+V(L_ACT1_6)*(0.011508)+V(L_ACT1_7)*(0.150744)+V(L_ACT1_8)*(-0.035876)+V(L_ACT1_9)*(0.090206)+V(L_ACT1_10)*(-0.219423)+V(L_ACT1_11)*(0.078821)+V(L_ACT1_12)*(-0.008443)+V(L_ACT1_13)*(0.096816)+V(L_ACT1_14)*(0.601903)+V(L_ACT1_15)*(-0.076234)+V(L_ACT1_16)*(0.020054)+V(L_ACT1_17)*(0.356409)+V(L_ACT1_18)*(0.239597)+V(L_ACT1_19)*(0.117298)+V(L_ACT1_20)*(0.250474)+V(L_ACT1_21)*(-0.162504)+V(L_ACT1_22)*(-0.146355)+V(L_ACT1_23)*(0.208444)+V(L_ACT1_24)*(0.069274)+V(L_ACT1_25)*(-0.328644)+V(L_ACT1_26)*(0.106269)+V(L_ACT1_27)*(0.215728)+V(L_ACT1_28)*(-0.056189)+V(L_ACT1_29)*(0.205561)+V(L_ACT1_30)*(0.075601)+V(L_ACT1_31)*(0.099760)+V(L_ACT1_32)*(-0.261296)+(0.110751))
B2_11 L2_11 0 V=(V(L_ACT1_1)*(0.309949)+V(L_ACT1_2)*(-0.162180)+V(L_ACT1_3)*(0.228457)+V(L_ACT1_4)*(-0.096997)+V(L_ACT1_5)*(0.122961)+V(L_ACT1_6)*(0.109062)+V(L_ACT1_7)*(0.171848)+V(L_ACT1_8)*(-0.230392)+V(L_ACT1_9)*(0.048734)+V(L_ACT1_10)*(0.053641)+V(L_ACT1_11)*(-0.015792)+V(L_ACT1_12)*(-0.058226)+V(L_ACT1_13)*(0.071371)+V(L_ACT1_14)*(0.610606)+V(L_ACT1_15)*(-0.207402)+V(L_ACT1_16)*(-0.010428)+V(L_ACT1_17)*(0.109880)+V(L_ACT1_18)*(0.209664)+V(L_ACT1_19)*(0.012627)+V(L_ACT1_20)*(0.059535)+V(L_ACT1_21)*(-0.072840)+V(L_ACT1_22)*(0.138066)+V(L_ACT1_23)*(0.260662)+V(L_ACT1_24)*(0.261743)+V(L_ACT1_25)*(-0.330832)+V(L_ACT1_26)*(0.013034)+V(L_ACT1_27)*(-0.114112)+V(L_ACT1_28)*(-0.085451)+V(L_ACT1_29)*(0.273516)+V(L_ACT1_30)*(0.214713)+V(L_ACT1_31)*(0.164430)+V(L_ACT1_32)*(-0.130172)+(0.119663))
B2_12 L2_12 0 V=(V(L_ACT1_1)*(0.010596)+V(L_ACT1_2)*(-0.110858)+V(L_ACT1_3)*(-0.114497)+V(L_ACT1_4)*(0.111964)+V(L_ACT1_5)*(-0.002387)+V(L_ACT1_6)*(0.005645)+V(L_ACT1_7)*(-0.025481)+V(L_ACT1_8)*(0.217957)+V(L_ACT1_9)*(-0.177741)+V(L_ACT1_10)*(0.072365)+V(L_ACT1_11)*(0.105958)+V(L_ACT1_12)*(-0.029978)+V(L_ACT1_13)*(-0.088669)+V(L_ACT1_14)*(0.008249)+V(L_ACT1_15)*(0.076127)+V(L_ACT1_16)*(0.242320)+V(L_ACT1_17)*(0.039053)+V(L_ACT1_18)*(0.153527)+V(L_ACT1_19)*(-0.205245)+V(L_ACT1_20)*(0.081468)+V(L_ACT1_21)*(0.226925)+V(L_ACT1_22)*(-0.008479)+V(L_ACT1_23)*(-0.002543)+V(L_ACT1_24)*(-0.008064)+V(L_ACT1_25)*(0.310357)+V(L_ACT1_26)*(-0.232547)+V(L_ACT1_27)*(-0.158433)+V(L_ACT1_28)*(0.029468)+V(L_ACT1_29)*(-0.059444)+V(L_ACT1_30)*(-0.007550)+V(L_ACT1_31)*(0.178270)+V(L_ACT1_32)*(-0.123805)+(-0.048995))
B2_13 L2_13 0 V=(V(L_ACT1_1)*(0.134092)+V(L_ACT1_2)*(0.087796)+V(L_ACT1_3)*(0.295101)+V(L_ACT1_4)*(0.124030)+V(L_ACT1_5)*(-0.132344)+V(L_ACT1_6)*(-0.082276)+V(L_ACT1_7)*(0.246635)+V(L_ACT1_8)*(-0.039712)+V(L_ACT1_9)*(-0.007380)+V(L_ACT1_10)*(-0.200282)+V(L_ACT1_11)*(0.054492)+V(L_ACT1_12)*(-0.232934)+V(L_ACT1_13)*(0.083631)+V(L_ACT1_14)*(0.468326)+V(L_ACT1_15)*(-0.234155)+V(L_ACT1_16)*(0.115297)+V(L_ACT1_17)*(0.345263)+V(L_ACT1_18)*(0.276643)+V(L_ACT1_19)*(0.160067)+V(L_ACT1_20)*(0.240269)+V(L_ACT1_21)*(-0.105025)+V(L_ACT1_22)*(-0.034951)+V(L_ACT1_23)*(0.023401)+V(L_ACT1_24)*(0.028002)+V(L_ACT1_25)*(-0.190796)+V(L_ACT1_26)*(0.135805)+V(L_ACT1_27)*(0.107159)+V(L_ACT1_28)*(-0.034210)+V(L_ACT1_29)*(0.171621)+V(L_ACT1_30)*(0.337872)+V(L_ACT1_31)*(0.258259)+V(L_ACT1_32)*(-0.338630)+(-0.001731))
B2_14 L2_14 0 V=(V(L_ACT1_1)*(0.059422)+V(L_ACT1_2)*(0.034844)+V(L_ACT1_3)*(-0.062256)+V(L_ACT1_4)*(0.178181)+V(L_ACT1_5)*(0.131550)+V(L_ACT1_6)*(0.112053)+V(L_ACT1_7)*(-0.256099)+V(L_ACT1_8)*(0.117453)+V(L_ACT1_9)*(-0.147315)+V(L_ACT1_10)*(0.226418)+V(L_ACT1_11)*(0.276498)+V(L_ACT1_12)*(0.253395)+V(L_ACT1_13)*(-0.026456)+V(L_ACT1_14)*(-0.306361)+V(L_ACT1_15)*(0.427803)+V(L_ACT1_16)*(0.258007)+V(L_ACT1_17)*(0.054458)+V(L_ACT1_18)*(-0.147644)+V(L_ACT1_19)*(0.004807)+V(L_ACT1_20)*(0.141269)+V(L_ACT1_21)*(0.182283)+V(L_ACT1_22)*(0.284964)+V(L_ACT1_23)*(-0.123553)+V(L_ACT1_24)*(0.043633)+V(L_ACT1_25)*(0.295727)+V(L_ACT1_26)*(0.019226)+V(L_ACT1_27)*(-0.191060)+V(L_ACT1_28)*(0.158470)+V(L_ACT1_29)*(-0.102420)+V(L_ACT1_30)*(-0.027182)+V(L_ACT1_31)*(-0.009284)+V(L_ACT1_32)*(0.343376)+(0.006347))
B2_15 L2_15 0 V=(V(L_ACT1_1)*(-0.216157)+V(L_ACT1_2)*(0.276330)+V(L_ACT1_3)*(-0.114371)+V(L_ACT1_4)*(0.230021)+V(L_ACT1_5)*(0.055292)+V(L_ACT1_6)*(0.264635)+V(L_ACT1_7)*(-0.185604)+V(L_ACT1_8)*(0.252258)+V(L_ACT1_9)*(-0.115521)+V(L_ACT1_10)*(0.276344)+V(L_ACT1_11)*(0.320175)+V(L_ACT1_12)*(0.298165)+V(L_ACT1_13)*(0.013566)+V(L_ACT1_14)*(-0.219854)+V(L_ACT1_15)*(0.199248)+V(L_ACT1_16)*(0.011059)+V(L_ACT1_17)*(0.000730)+V(L_ACT1_18)*(-0.046944)+V(L_ACT1_19)*(-0.125729)+V(L_ACT1_20)*(-0.064530)+V(L_ACT1_21)*(0.106193)+V(L_ACT1_22)*(0.226904)+V(L_ACT1_23)*(-0.050836)+V(L_ACT1_24)*(-0.048370)+V(L_ACT1_25)*(0.330560)+V(L_ACT1_26)*(0.202069)+V(L_ACT1_27)*(-0.071016)+V(L_ACT1_28)*(0.032947)+V(L_ACT1_29)*(-0.197642)+V(L_ACT1_30)*(0.018380)+V(L_ACT1_31)*(-0.038955)+V(L_ACT1_32)*(0.037338)+(0.215912))
B2_16 L2_16 0 V=(V(L_ACT1_1)*(-0.124534)+V(L_ACT1_2)*(0.253901)+V(L_ACT1_3)*(-0.072672)+V(L_ACT1_4)*(0.330902)+V(L_ACT1_5)*(0.263208)+V(L_ACT1_6)*(0.025336)+V(L_ACT1_7)*(-0.193564)+V(L_ACT1_8)*(-0.012778)+V(L_ACT1_9)*(-0.138821)+V(L_ACT1_10)*(0.054119)+V(L_ACT1_11)*(0.251129)+V(L_ACT1_12)*(0.323882)+V(L_ACT1_13)*(0.199566)+V(L_ACT1_14)*(-0.179808)+V(L_ACT1_15)*(0.411822)+V(L_ACT1_16)*(0.089335)+V(L_ACT1_17)*(0.044238)+V(L_ACT1_18)*(0.057469)+V(L_ACT1_19)*(-0.079691)+V(L_ACT1_20)*(-0.072588)+V(L_ACT1_21)*(0.229761)+V(L_ACT1_22)*(0.164191)+V(L_ACT1_23)*(0.125499)+V(L_ACT1_24)*(-0.183389)+V(L_ACT1_25)*(0.343048)+V(L_ACT1_26)*(0.010773)+V(L_ACT1_27)*(0.114018)+V(L_ACT1_28)*(0.187328)+V(L_ACT1_29)*(-0.295944)+V(L_ACT1_30)*(-0.131083)+V(L_ACT1_31)*(-0.199985)+V(L_ACT1_32)*(0.128688)+(0.034075))
* ACTIVATION LAYER 2: RELU
B_ACT2_1 L_ACT2_1 0 V=(IF(V(L2_1)>0,V(L2_1),0))
B_ACT2_2 L_ACT2_2 0 V=(IF(V(L2_2)>0,V(L2_2),0))
B_ACT2_3 L_ACT2_3 0 V=(IF(V(L2_3)>0,V(L2_3),0))
B_ACT2_4 L_ACT2_4 0 V=(IF(V(L2_4)>0,V(L2_4),0))
B_ACT2_5 L_ACT2_5 0 V=(IF(V(L2_5)>0,V(L2_5),0))
B_ACT2_6 L_ACT2_6 0 V=(IF(V(L2_6)>0,V(L2_6),0))
B_ACT2_7 L_ACT2_7 0 V=(IF(V(L2_7)>0,V(L2_7),0))
B_ACT2_8 L_ACT2_8 0 V=(IF(V(L2_8)>0,V(L2_8),0))
B_ACT2_9 L_ACT2_9 0 V=(IF(V(L2_9)>0,V(L2_9),0))
B_ACT2_10 L_ACT2_10 0 V=(IF(V(L2_10)>0,V(L2_10),0))
B_ACT2_11 L_ACT2_11 0 V=(IF(V(L2_11)>0,V(L2_11),0))
B_ACT2_12 L_ACT2_12 0 V=(IF(V(L2_12)>0,V(L2_12),0))
B_ACT2_13 L_ACT2_13 0 V=(IF(V(L2_13)>0,V(L2_13),0))
B_ACT2_14 L_ACT2_14 0 V=(IF(V(L2_14)>0,V(L2_14),0))
B_ACT2_15 L_ACT2_15 0 V=(IF(V(L2_15)>0,V(L2_15),0))
B_ACT2_16 L_ACT2_16 0 V=(IF(V(L2_16)>0,V(L2_16),0))
* LAYER 3: LINEAR
B3_1 L3_1 0 V=(V(L_ACT2_1)*(0.265448)+V(L_ACT2_2)*(0.306892)+V(L_ACT2_3)*(-0.132897)+V(L_ACT2_4)*(-0.232571)+V(L_ACT2_5)*(-0.264658)+V(L_ACT2_6)*(-0.321262)+V(L_ACT2_7)*(0.040762)+V(L_ACT2_8)*(-0.387965)+V(L_ACT2_9)*(-0.839529)+V(L_ACT2_10)*(-0.346777)+V(L_ACT2_11)*(-0.365063)+V(L_ACT2_12)*(0.188376)+V(L_ACT2_13)*(-0.249895)+V(L_ACT2_14)*(0.340903)+V(L_ACT2_15)*(0.372237)+V(L_ACT2_16)*(0.291442)+(0.008520))
* ACTIVATION LAYER 3: SIGMOID
B_ACT3_1 L_ACT3_1 0 V=(1/(1+EXP(-V(L3_1))))
* Connect final internal node L_ACT3_1 to external output NNOUT1
B_OUT NNOUT1 0 V=V(L_ACT3_1)
.ENDS ActorSubckt