.SUBCKT ActorSubckt NNIN1 NNIN2 NNIN3 NNIN4 NNIN5 NNIN6 NNIN7 NNIN8 NNIN9 NNIN10 NNIN11 NNIN12 NNIN13 NNIN14 NNIN15 NNIN16 NNIN17 NNIN18 NNIN19 NNOUT1

* LAYER 1: LINEAR
B1_1 L1_1 0 V=(V(NNIN1)*(-0.081883)+V(NNIN2)*(0.114159)+V(NNIN3)*(-0.114844)+V(NNIN4)*(-0.003784)+V(NNIN5)*(-0.220726)+V(NNIN6)*(0.554409)+V(NNIN7)*(0.888378)+V(NNIN8)*(0.647330)+V(NNIN9)*(0.484143)+V(NNIN10)*(0.572619)+V(NNIN11)*(-0.459769)+V(NNIN12)*(-0.059756)+V(NNIN13)*(0.067945)+V(NNIN14)*(0.050554)+V(NNIN15)*(-0.103654)+V(NNIN16)*(0.234317)+V(NNIN17)*(0.013964)+V(NNIN18)*(-0.335066)+V(NNIN19)*(-0.150129)+(0.135601))
B1_2 L1_2 0 V=(V(NNIN1)*(0.045873)+V(NNIN2)*(0.125584)+V(NNIN3)*(-0.208204)+V(NNIN4)*(0.020089)+V(NNIN5)*(0.054018)+V(NNIN6)*(1.271392)+V(NNIN7)*(0.952228)+V(NNIN8)*(1.068899)+V(NNIN9)*(0.739231)+V(NNIN10)*(0.809097)+V(NNIN11)*(-0.066302)+V(NNIN12)*(-0.235378)+V(NNIN13)*(0.183376)+V(NNIN14)*(-0.168572)+V(NNIN15)*(-0.027914)+V(NNIN16)*(0.094062)+V(NNIN17)*(0.039873)+V(NNIN18)*(-0.188022)+V(NNIN19)*(-0.219615)+(0.211062))
B1_3 L1_3 0 V=(V(NNIN1)*(0.149369)+V(NNIN2)*(0.138050)+V(NNIN3)*(0.265011)+V(NNIN4)*(0.464842)+V(NNIN5)*(0.130309)+V(NNIN6)*(-0.107434)+V(NNIN7)*(0.299606)+V(NNIN8)*(0.378879)+V(NNIN9)*(0.497992)+V(NNIN10)*(0.483665)+V(NNIN11)*(-0.293513)+V(NNIN12)*(-0.229792)+V(NNIN13)*(0.136715)+V(NNIN14)*(0.178597)+V(NNIN15)*(0.000901)+V(NNIN16)*(0.413134)+V(NNIN17)*(0.318047)+V(NNIN18)*(-0.092324)+V(NNIN19)*(0.483794)+(0.385313))
B1_4 L1_4 0 V=(V(NNIN1)*(0.471027)+V(NNIN2)*(0.493654)+V(NNIN3)*(0.383780)+V(NNIN4)*(0.179059)+V(NNIN5)*(0.312597)+V(NNIN6)*(-1.367919)+V(NNIN7)*(-1.142584)+V(NNIN8)*(-0.636932)+V(NNIN9)*(-0.848743)+V(NNIN10)*(-0.469395)+V(NNIN11)*(0.177014)+V(NNIN12)*(0.101652)+V(NNIN13)*(0.377521)+V(NNIN14)*(0.268547)+V(NNIN15)*(0.111512)+V(NNIN16)*(0.021150)+V(NNIN17)*(0.372189)+V(NNIN18)*(0.308311)+V(NNIN19)*(-0.098095)+(0.115243))
B1_5 L1_5 0 V=(V(NNIN1)*(-0.133404)+V(NNIN2)*(0.120691)+V(NNIN3)*(0.185744)+V(NNIN4)*(0.043194)+V(NNIN5)*(-0.099209)+V(NNIN6)*(1.124997)+V(NNIN7)*(0.894499)+V(NNIN8)*(0.883393)+V(NNIN9)*(0.537814)+V(NNIN10)*(0.750964)+V(NNIN11)*(-0.005247)+V(NNIN12)*(-0.094524)+V(NNIN13)*(0.166112)+V(NNIN14)*(-0.178213)+V(NNIN15)*(0.054819)+V(NNIN16)*(0.096671)+V(NNIN17)*(0.169945)+V(NNIN18)*(-0.462987)+V(NNIN19)*(-0.260393)+(0.082323))
B1_6 L1_6 0 V=(V(NNIN1)*(-0.053956)+V(NNIN2)*(0.112541)+V(NNIN3)*(0.211472)+V(NNIN4)*(0.024348)+V(NNIN5)*(-0.155449)+V(NNIN6)*(0.754220)+V(NNIN7)*(0.897549)+V(NNIN8)*(0.439327)+V(NNIN9)*(0.335331)+V(NNIN10)*(0.219271)+V(NNIN11)*(-0.111796)+V(NNIN12)*(-0.026166)+V(NNIN13)*(0.179855)+V(NNIN14)*(0.074894)+V(NNIN15)*(-0.024856)+V(NNIN16)*(-0.110169)+V(NNIN17)*(-0.159897)+V(NNIN18)*(-0.054317)+V(NNIN19)*(-0.268255)+(0.174551))
B1_7 L1_7 0 V=(V(NNIN1)*(0.192143)+V(NNIN2)*(0.050427)+V(NNIN3)*(0.118073)+V(NNIN4)*(0.086833)+V(NNIN5)*(0.200571)+V(NNIN6)*(0.100426)+V(NNIN7)*(0.283035)+V(NNIN8)*(0.434067)+V(NNIN9)*(0.664454)+V(NNIN10)*(0.758876)+V(NNIN11)*(-0.107339)+V(NNIN12)*(-0.005962)+V(NNIN13)*(-0.096237)+V(NNIN14)*(0.083527)+V(NNIN15)*(-0.172650)+V(NNIN16)*(0.295426)+V(NNIN17)*(0.054614)+V(NNIN18)*(-0.060552)+V(NNIN19)*(0.515685)+(-0.060762))
B1_8 L1_8 0 V=(V(NNIN1)*(-0.163092)+V(NNIN2)*(-0.054575)+V(NNIN3)*(0.225032)+V(NNIN4)*(0.182834)+V(NNIN5)*(-0.123198)+V(NNIN6)*(0.433268)+V(NNIN7)*(0.388151)+V(NNIN8)*(0.147244)+V(NNIN9)*(0.207207)+V(NNIN10)*(0.397329)+V(NNIN11)*(-0.277531)+V(NNIN12)*(-0.146286)+V(NNIN13)*(0.034734)+V(NNIN14)*(-0.065237)+V(NNIN15)*(-0.178188)+V(NNIN16)*(-0.035670)+V(NNIN17)*(-0.121531)+V(NNIN18)*(-0.288636)+V(NNIN19)*(-0.173791)+(0.211308))
B1_9 L1_9 0 V=(V(NNIN1)*(0.099054)+V(NNIN2)*(0.105562)+V(NNIN3)*(0.250438)+V(NNIN4)*(0.232583)+V(NNIN5)*(0.131412)+V(NNIN6)*(1.419782)+V(NNIN7)*(1.334751)+V(NNIN8)*(1.072032)+V(NNIN9)*(0.792049)+V(NNIN10)*(0.856944)+V(NNIN11)*(-0.025063)+V(NNIN12)*(-0.093967)+V(NNIN13)*(0.222650)+V(NNIN14)*(0.025789)+V(NNIN15)*(0.050284)+V(NNIN16)*(-0.087910)+V(NNIN17)*(0.076733)+V(NNIN18)*(-0.026494)+V(NNIN19)*(0.106920)+(-0.044526))
B1_10 L1_10 0 V=(V(NNIN1)*(0.196516)+V(NNIN2)*(-0.177348)+V(NNIN3)*(0.013673)+V(NNIN4)*(-0.003288)+V(NNIN5)*(0.163913)+V(NNIN6)*(0.520811)+V(NNIN7)*(0.406404)+V(NNIN8)*(0.216430)+V(NNIN9)*(0.354627)+V(NNIN10)*(0.304147)+V(NNIN11)*(-0.243726)+V(NNIN12)*(-0.399817)+V(NNIN13)*(-0.198544)+V(NNIN14)*(-0.199174)+V(NNIN15)*(0.006368)+V(NNIN16)*(-0.107476)+V(NNIN17)*(-0.008578)+V(NNIN18)*(-0.093663)+V(NNIN19)*(-0.214622)+(-0.096968))
B1_11 L1_11 0 V=(V(NNIN1)*(0.223980)+V(NNIN2)*(0.242275)+V(NNIN3)*(0.183918)+V(NNIN4)*(-0.149336)+V(NNIN5)*(0.217929)+V(NNIN6)*(1.269647)+V(NNIN7)*(1.558603)+V(NNIN8)*(1.267537)+V(NNIN9)*(1.125368)+V(NNIN10)*(0.853545)+V(NNIN11)*(0.019920)+V(NNIN12)*(0.056659)+V(NNIN13)*(-0.047314)+V(NNIN14)*(0.103187)+V(NNIN15)*(0.127741)+V(NNIN16)*(0.085507)+V(NNIN17)*(-0.010079)+V(NNIN18)*(-0.335893)+V(NNIN19)*(0.066647)+(0.016486))
B1_12 L1_12 0 V=(V(NNIN1)*(0.295066)+V(NNIN2)*(0.042659)+V(NNIN3)*(0.245036)+V(NNIN4)*(0.300964)+V(NNIN5)*(0.178776)+V(NNIN6)*(1.547561)+V(NNIN7)*(1.323607)+V(NNIN8)*(1.233251)+V(NNIN9)*(0.960124)+V(NNIN10)*(0.619817)+V(NNIN11)*(-0.149922)+V(NNIN12)*(0.041506)+V(NNIN13)*(0.098996)+V(NNIN14)*(0.193060)+V(NNIN15)*(0.077638)+V(NNIN16)*(0.144089)+V(NNIN17)*(0.084380)+V(NNIN18)*(-0.128393)+V(NNIN19)*(0.137086)+(-0.030504))
B1_13 L1_13 0 V=(V(NNIN1)*(0.072657)+V(NNIN2)*(-0.149275)+V(NNIN3)*(0.235502)+V(NNIN4)*(-0.075186)+V(NNIN5)*(0.118072)+V(NNIN6)*(1.284368)+V(NNIN7)*(1.332320)+V(NNIN8)*(0.763117)+V(NNIN9)*(0.743411)+V(NNIN10)*(0.720260)+V(NNIN11)*(0.094277)+V(NNIN12)*(0.127424)+V(NNIN13)*(-0.090147)+V(NNIN14)*(0.086305)+V(NNIN15)*(0.095315)+V(NNIN16)*(0.348387)+V(NNIN17)*(-0.132329)+V(NNIN18)*(-0.097072)+V(NNIN19)*(0.173178)+(0.157464))
B1_14 L1_14 0 V=(V(NNIN1)*(0.051299)+V(NNIN2)*(0.140018)+V(NNIN3)*(0.051154)+V(NNIN4)*(0.199979)+V(NNIN5)*(0.246674)+V(NNIN6)*(-1.057889)+V(NNIN7)*(-0.913913)+V(NNIN8)*(-0.827317)+V(NNIN9)*(-0.585034)+V(NNIN10)*(-0.583938)+V(NNIN11)*(0.496790)+V(NNIN12)*(0.136940)+V(NNIN13)*(0.090939)+V(NNIN14)*(0.254816)+V(NNIN15)*(0.360502)+V(NNIN16)*(0.233435)+V(NNIN17)*(0.529413)+V(NNIN18)*(0.108245)+V(NNIN19)*(-0.125173)+(0.232797))
B1_15 L1_15 0 V=(V(NNIN1)*(-0.146793)+V(NNIN2)*(-0.054101)+V(NNIN3)*(-0.230971)+V(NNIN4)*(0.048500)+V(NNIN5)*(-0.041680)+V(NNIN6)*(0.488761)+V(NNIN7)*(0.592588)+V(NNIN8)*(0.368199)+V(NNIN9)*(0.111051)+V(NNIN10)*(0.006055)+V(NNIN11)*(0.113902)+V(NNIN12)*(0.060366)+V(NNIN13)*(-0.135928)+V(NNIN14)*(0.116022)+V(NNIN15)*(-0.034498)+V(NNIN16)*(0.034579)+V(NNIN17)*(-0.236059)+V(NNIN18)*(0.213653)+V(NNIN19)*(0.104576)+(0.335714))
B1_16 L1_16 0 V=(V(NNIN1)*(-0.135162)+V(NNIN2)*(0.216582)+V(NNIN3)*(-0.088135)+V(NNIN4)*(-0.209198)+V(NNIN5)*(-0.164795)+V(NNIN6)*(1.067261)+V(NNIN7)*(0.896933)+V(NNIN8)*(0.354753)+V(NNIN9)*(0.275107)+V(NNIN10)*(0.243085)+V(NNIN11)*(0.225068)+V(NNIN12)*(0.081078)+V(NNIN13)*(0.158568)+V(NNIN14)*(-0.136014)+V(NNIN15)*(0.083503)+V(NNIN16)*(0.234511)+V(NNIN17)*(-0.130206)+V(NNIN18)*(-0.155485)+V(NNIN19)*(0.310572)+(0.200322))
B1_17 L1_17 0 V=(V(NNIN1)*(0.168146)+V(NNIN2)*(0.120432)+V(NNIN3)*(0.088657)+V(NNIN4)*(-0.109601)+V(NNIN5)*(-0.126960)+V(NNIN6)*(1.471464)+V(NNIN7)*(1.157866)+V(NNIN8)*(0.895560)+V(NNIN9)*(1.008124)+V(NNIN10)*(0.516861)+V(NNIN11)*(-0.148696)+V(NNIN12)*(-0.050918)+V(NNIN13)*(0.269480)+V(NNIN14)*(0.295581)+V(NNIN15)*(0.164050)+V(NNIN16)*(0.372143)+V(NNIN17)*(-0.110592)+V(NNIN18)*(-0.007872)+V(NNIN19)*(0.103288)+(0.117283))
B1_18 L1_18 0 V=(V(NNIN1)*(-0.137531)+V(NNIN2)*(-0.065116)+V(NNIN3)*(0.199867)+V(NNIN4)*(-0.165688)+V(NNIN5)*(-0.007106)+V(NNIN6)*(1.090399)+V(NNIN7)*(0.853203)+V(NNIN8)*(0.548124)+V(NNIN9)*(0.677393)+V(NNIN10)*(0.347595)+V(NNIN11)*(-0.164425)+V(NNIN12)*(-0.024726)+V(NNIN13)*(0.287603)+V(NNIN14)*(0.066988)+V(NNIN15)*(-0.112091)+V(NNIN16)*(0.357907)+V(NNIN17)*(-0.071200)+V(NNIN18)*(-0.047337)+V(NNIN19)*(0.332619)+(0.237442))
B1_19 L1_19 0 V=(V(NNIN1)*(-0.020336)+V(NNIN2)*(0.131329)+V(NNIN3)*(-0.024226)+V(NNIN4)*(-0.049479)+V(NNIN5)*(0.230264)+V(NNIN6)*(-1.049157)+V(NNIN7)*(-1.148427)+V(NNIN8)*(-0.986916)+V(NNIN9)*(-0.786430)+V(NNIN10)*(-0.797414)+V(NNIN11)*(0.187426)+V(NNIN12)*(0.316625)+V(NNIN13)*(0.004699)+V(NNIN14)*(0.061845)+V(NNIN15)*(-0.019200)+V(NNIN16)*(0.228648)+V(NNIN17)*(0.055886)+V(NNIN18)*(0.047172)+V(NNIN19)*(0.015677)+(0.169495))
B1_20 L1_20 0 V=(V(NNIN1)*(0.064444)+V(NNIN2)*(0.086628)+V(NNIN3)*(0.340863)+V(NNIN4)*(0.271383)+V(NNIN5)*(0.024275)+V(NNIN6)*(1.448041)+V(NNIN7)*(0.990035)+V(NNIN8)*(1.094688)+V(NNIN9)*(0.871008)+V(NNIN10)*(0.743309)+V(NNIN11)*(-0.239437)+V(NNIN12)*(0.170665)+V(NNIN13)*(0.172871)+V(NNIN14)*(0.226915)+V(NNIN15)*(0.011169)+V(NNIN16)*(0.231634)+V(NNIN17)*(0.074806)+V(NNIN18)*(0.019701)+V(NNIN19)*(0.239765)+(0.129910))
B1_21 L1_21 0 V=(V(NNIN1)*(0.494271)+V(NNIN2)*(0.472576)+V(NNIN3)*(0.114557)+V(NNIN4)*(0.153216)+V(NNIN5)*(0.188356)+V(NNIN6)*(-1.198660)+V(NNIN7)*(-0.799918)+V(NNIN8)*(-0.751133)+V(NNIN9)*(-0.289535)+V(NNIN10)*(-0.159749)+V(NNIN11)*(0.274178)+V(NNIN12)*(-0.007901)+V(NNIN13)*(0.001649)+V(NNIN14)*(0.185511)+V(NNIN15)*(0.140620)+V(NNIN16)*(0.434317)+V(NNIN17)*(0.209711)+V(NNIN18)*(-0.157057)+V(NNIN19)*(0.105206)+(0.268843))
B1_22 L1_22 0 V=(V(NNIN1)*(-0.027964)+V(NNIN2)*(-0.047221)+V(NNIN3)*(-0.014736)+V(NNIN4)*(-0.025956)+V(NNIN5)*(0.141629)+V(NNIN6)*(-0.018216)+V(NNIN7)*(-0.348631)+V(NNIN8)*(-0.043260)+V(NNIN9)*(-0.058875)+V(NNIN10)*(-0.171567)+V(NNIN11)*(0.220554)+V(NNIN12)*(0.048626)+V(NNIN13)*(0.077315)+V(NNIN14)*(0.012426)+V(NNIN15)*(0.164056)+V(NNIN16)*(-0.251510)+V(NNIN17)*(-0.143118)+V(NNIN18)*(0.257375)+V(NNIN19)*(0.179126)+(-0.219540))
B1_23 L1_23 0 V=(V(NNIN1)*(0.418787)+V(NNIN2)*(0.399322)+V(NNIN3)*(0.058046)+V(NNIN4)*(0.052087)+V(NNIN5)*(0.242430)+V(NNIN6)*(-1.064929)+V(NNIN7)*(-0.873722)+V(NNIN8)*(-0.786051)+V(NNIN9)*(-0.655699)+V(NNIN10)*(-0.584664)+V(NNIN11)*(0.401554)+V(NNIN12)*(0.255110)+V(NNIN13)*(0.022028)+V(NNIN14)*(0.244750)+V(NNIN15)*(0.335227)+V(NNIN16)*(0.006695)+V(NNIN17)*(0.193609)+V(NNIN18)*(0.405618)+V(NNIN19)*(0.075484)+(0.177944))
B1_24 L1_24 0 V=(V(NNIN1)*(-0.064032)+V(NNIN2)*(0.051099)+V(NNIN3)*(0.238548)+V(NNIN4)*(0.131725)+V(NNIN5)*(0.096239)+V(NNIN6)*(1.070744)+V(NNIN7)*(0.803035)+V(NNIN8)*(0.646051)+V(NNIN9)*(0.567717)+V(NNIN10)*(0.789889)+V(NNIN11)*(-0.135921)+V(NNIN12)*(-0.099128)+V(NNIN13)*(-0.180532)+V(NNIN14)*(-0.002247)+V(NNIN15)*(-0.261922)+V(NNIN16)*(0.205776)+V(NNIN17)*(-0.083250)+V(NNIN18)*(0.049192)+V(NNIN19)*(0.067779)+(0.162253))
B1_25 L1_25 0 V=(V(NNIN1)*(0.099275)+V(NNIN2)*(0.109928)+V(NNIN3)*(0.141371)+V(NNIN4)*(0.092020)+V(NNIN5)*(-0.045300)+V(NNIN6)*(1.689185)+V(NNIN7)*(1.433238)+V(NNIN8)*(1.235423)+V(NNIN9)*(0.718947)+V(NNIN10)*(0.959373)+V(NNIN11)*(-0.299346)+V(NNIN12)*(0.184953)+V(NNIN13)*(0.001441)+V(NNIN14)*(0.210945)+V(NNIN15)*(0.240273)+V(NNIN16)*(0.146265)+V(NNIN17)*(0.157559)+V(NNIN18)*(-0.315382)+V(NNIN19)*(0.100169)+(0.206008))
B1_26 L1_26 0 V=(V(NNIN1)*(-0.044860)+V(NNIN2)*(-0.282395)+V(NNIN3)*(0.036303)+V(NNIN4)*(-0.287527)+V(NNIN5)*(-0.171612)+V(NNIN6)*(0.855056)+V(NNIN7)*(0.637429)+V(NNIN8)*(0.699709)+V(NNIN9)*(0.692334)+V(NNIN10)*(0.400547)+V(NNIN11)*(-0.051271)+V(NNIN12)*(-0.094027)+V(NNIN13)*(0.309616)+V(NNIN14)*(-0.015566)+V(NNIN15)*(0.218615)+V(NNIN16)*(0.214510)+V(NNIN17)*(-0.305383)+V(NNIN18)*(-0.268216)+V(NNIN19)*(0.223523)+(0.009766))
B1_27 L1_27 0 V=(V(NNIN1)*(0.171787)+V(NNIN2)*(0.075877)+V(NNIN3)*(0.105307)+V(NNIN4)*(-0.200284)+V(NNIN5)*(-0.230207)+V(NNIN6)*(0.772318)+V(NNIN7)*(0.824226)+V(NNIN8)*(1.106020)+V(NNIN9)*(0.868928)+V(NNIN10)*(0.633880)+V(NNIN11)*(-0.515250)+V(NNIN12)*(-0.340076)+V(NNIN13)*(0.023184)+V(NNIN14)*(0.077163)+V(NNIN15)*(0.116224)+V(NNIN16)*(0.275362)+V(NNIN17)*(0.069358)+V(NNIN18)*(-0.387206)+V(NNIN19)*(-0.249531)+(0.072412))
B1_28 L1_28 0 V=(V(NNIN1)*(0.011354)+V(NNIN2)*(0.072375)+V(NNIN3)*(-0.068642)+V(NNIN4)*(-0.132677)+V(NNIN5)*(-0.028126)+V(NNIN6)*(0.876275)+V(NNIN7)*(1.032294)+V(NNIN8)*(0.938567)+V(NNIN9)*(0.716182)+V(NNIN10)*(0.534016)+V(NNIN11)*(0.229396)+V(NNIN12)*(0.063659)+V(NNIN13)*(0.121937)+V(NNIN14)*(0.016707)+V(NNIN15)*(0.128815)+V(NNIN16)*(0.138843)+V(NNIN17)*(-0.155320)+V(NNIN18)*(-0.023300)+V(NNIN19)*(0.171101)+(0.118471))
B1_29 L1_29 0 V=(V(NNIN1)*(0.166086)+V(NNIN2)*(0.174905)+V(NNIN3)*(-0.068242)+V(NNIN4)*(0.253415)+V(NNIN5)*(-0.145533)+V(NNIN6)*(1.069588)+V(NNIN7)*(0.871662)+V(NNIN8)*(0.786027)+V(NNIN9)*(0.804224)+V(NNIN10)*(0.761472)+V(NNIN11)*(0.254364)+V(NNIN12)*(-0.130097)+V(NNIN13)*(0.030296)+V(NNIN14)*(-0.003406)+V(NNIN15)*(0.042538)+V(NNIN16)*(-0.081356)+V(NNIN17)*(0.001369)+V(NNIN18)*(-0.029888)+V(NNIN19)*(-0.111366)+(-0.092520))
B1_30 L1_30 0 V=(V(NNIN1)*(-0.218413)+V(NNIN2)*(-0.174896)+V(NNIN3)*(-0.030906)+V(NNIN4)*(0.090531)+V(NNIN5)*(-0.090407)+V(NNIN6)*(0.858558)+V(NNIN7)*(0.754224)+V(NNIN8)*(0.775548)+V(NNIN9)*(0.728459)+V(NNIN10)*(0.564347)+V(NNIN11)*(-0.387124)+V(NNIN12)*(-0.132312)+V(NNIN13)*(-0.145801)+V(NNIN14)*(0.049752)+V(NNIN15)*(0.057154)+V(NNIN16)*(0.310976)+V(NNIN17)*(0.127346)+V(NNIN18)*(-0.324598)+V(NNIN19)*(-0.219758)+(0.138346))
B1_31 L1_31 0 V=(V(NNIN1)*(0.186887)+V(NNIN2)*(0.054634)+V(NNIN3)*(0.246465)+V(NNIN4)*(0.215738)+V(NNIN5)*(-0.196691)+V(NNIN6)*(1.508730)+V(NNIN7)*(1.287984)+V(NNIN8)*(1.180752)+V(NNIN9)*(0.724459)+V(NNIN10)*(0.738371)+V(NNIN11)*(-0.048208)+V(NNIN12)*(0.237430)+V(NNIN13)*(0.291237)+V(NNIN14)*(0.158080)+V(NNIN15)*(0.120847)+V(NNIN16)*(0.275535)+V(NNIN17)*(0.095608)+V(NNIN18)*(-0.147073)+V(NNIN19)*(0.069937)+(-0.104522))
B1_32 L1_32 0 V=(V(NNIN1)*(0.149330)+V(NNIN2)*(-0.129621)+V(NNIN3)*(-0.194795)+V(NNIN4)*(-0.103434)+V(NNIN5)*(-0.044088)+V(NNIN6)*(0.395292)+V(NNIN7)*(0.633267)+V(NNIN8)*(0.416864)+V(NNIN9)*(0.206050)+V(NNIN10)*(0.109418)+V(NNIN11)*(0.158132)+V(NNIN12)*(0.126271)+V(NNIN13)*(-0.103986)+V(NNIN14)*(0.171122)+V(NNIN15)*(0.089221)+V(NNIN16)*(-0.124691)+V(NNIN17)*(0.124234)+V(NNIN18)*(-0.121642)+V(NNIN19)*(-0.136011)+(-0.230807))
* ACTIVATION LAYER 1: RELU
B_ACT1_1 L_ACT1_1 0 V=(IF(V(L1_1)>0,V(L1_1),0))
B_ACT1_2 L_ACT1_2 0 V=(IF(V(L1_2)>0,V(L1_2),0))
B_ACT1_3 L_ACT1_3 0 V=(IF(V(L1_3)>0,V(L1_3),0))
B_ACT1_4 L_ACT1_4 0 V=(IF(V(L1_4)>0,V(L1_4),0))
B_ACT1_5 L_ACT1_5 0 V=(IF(V(L1_5)>0,V(L1_5),0))
B_ACT1_6 L_ACT1_6 0 V=(IF(V(L1_6)>0,V(L1_6),0))
B_ACT1_7 L_ACT1_7 0 V=(IF(V(L1_7)>0,V(L1_7),0))
B_ACT1_8 L_ACT1_8 0 V=(IF(V(L1_8)>0,V(L1_8),0))
B_ACT1_9 L_ACT1_9 0 V=(IF(V(L1_9)>0,V(L1_9),0))
B_ACT1_10 L_ACT1_10 0 V=(IF(V(L1_10)>0,V(L1_10),0))
B_ACT1_11 L_ACT1_11 0 V=(IF(V(L1_11)>0,V(L1_11),0))
B_ACT1_12 L_ACT1_12 0 V=(IF(V(L1_12)>0,V(L1_12),0))
B_ACT1_13 L_ACT1_13 0 V=(IF(V(L1_13)>0,V(L1_13),0))
B_ACT1_14 L_ACT1_14 0 V=(IF(V(L1_14)>0,V(L1_14),0))
B_ACT1_15 L_ACT1_15 0 V=(IF(V(L1_15)>0,V(L1_15),0))
B_ACT1_16 L_ACT1_16 0 V=(IF(V(L1_16)>0,V(L1_16),0))
B_ACT1_17 L_ACT1_17 0 V=(IF(V(L1_17)>0,V(L1_17),0))
B_ACT1_18 L_ACT1_18 0 V=(IF(V(L1_18)>0,V(L1_18),0))
B_ACT1_19 L_ACT1_19 0 V=(IF(V(L1_19)>0,V(L1_19),0))
B_ACT1_20 L_ACT1_20 0 V=(IF(V(L1_20)>0,V(L1_20),0))
B_ACT1_21 L_ACT1_21 0 V=(IF(V(L1_21)>0,V(L1_21),0))
B_ACT1_22 L_ACT1_22 0 V=(IF(V(L1_22)>0,V(L1_22),0))
B_ACT1_23 L_ACT1_23 0 V=(IF(V(L1_23)>0,V(L1_23),0))
B_ACT1_24 L_ACT1_24 0 V=(IF(V(L1_24)>0,V(L1_24),0))
B_ACT1_25 L_ACT1_25 0 V=(IF(V(L1_25)>0,V(L1_25),0))
B_ACT1_26 L_ACT1_26 0 V=(IF(V(L1_26)>0,V(L1_26),0))
B_ACT1_27 L_ACT1_27 0 V=(IF(V(L1_27)>0,V(L1_27),0))
B_ACT1_28 L_ACT1_28 0 V=(IF(V(L1_28)>0,V(L1_28),0))
B_ACT1_29 L_ACT1_29 0 V=(IF(V(L1_29)>0,V(L1_29),0))
B_ACT1_30 L_ACT1_30 0 V=(IF(V(L1_30)>0,V(L1_30),0))
B_ACT1_31 L_ACT1_31 0 V=(IF(V(L1_31)>0,V(L1_31),0))
B_ACT1_32 L_ACT1_32 0 V=(IF(V(L1_32)>0,V(L1_32),0))
* LAYER 2: LINEAR
B2_1 L2_1 0 V=(V(L_ACT1_1)*(-0.546027)+V(L_ACT1_2)*(0.124211)+V(L_ACT1_3)*(0.225769)+V(L_ACT1_4)*(0.165019)+V(L_ACT1_5)*(-0.218020)+V(L_ACT1_6)*(-0.200137)+V(L_ACT1_7)*(0.244328)+V(L_ACT1_8)*(-0.214161)+V(L_ACT1_9)*(-0.043683)+V(L_ACT1_10)*(-0.096297)+V(L_ACT1_11)*(-0.052127)+V(L_ACT1_12)*(-0.025486)+V(L_ACT1_13)*(0.190549)+V(L_ACT1_14)*(0.028884)+V(L_ACT1_15)*(-0.122070)+V(L_ACT1_16)*(-0.333304)+V(L_ACT1_17)*(0.014945)+V(L_ACT1_18)*(-0.102772)+V(L_ACT1_19)*(0.153875)+V(L_ACT1_20)*(0.080907)+V(L_ACT1_21)*(0.148284)+V(L_ACT1_22)*(-0.161459)+V(L_ACT1_23)*(0.183307)+V(L_ACT1_24)*(-0.181239)+V(L_ACT1_25)*(-0.052706)+V(L_ACT1_26)*(-0.172860)+V(L_ACT1_27)*(0.004540)+V(L_ACT1_28)*(-0.229345)+V(L_ACT1_29)*(-0.275597)+V(L_ACT1_30)*(-0.342783)+V(L_ACT1_31)*(0.015583)+V(L_ACT1_32)*(-0.287247)+(0.246171))
B2_2 L2_2 0 V=(V(L_ACT1_1)*(0.465762)+V(L_ACT1_2)*(0.015132)+V(L_ACT1_3)*(0.225099)+V(L_ACT1_4)*(0.116009)+V(L_ACT1_5)*(0.228092)+V(L_ACT1_6)*(0.318770)+V(L_ACT1_7)*(0.159951)+V(L_ACT1_8)*(0.281214)+V(L_ACT1_9)*(0.332998)+V(L_ACT1_10)*(0.040798)+V(L_ACT1_11)*(0.179182)+V(L_ACT1_12)*(0.092663)+V(L_ACT1_13)*(0.319630)+V(L_ACT1_14)*(-0.149987)+V(L_ACT1_15)*(0.184643)+V(L_ACT1_16)*(0.334905)+V(L_ACT1_17)*(0.414173)+V(L_ACT1_18)*(0.330736)+V(L_ACT1_19)*(-0.082004)+V(L_ACT1_20)*(-0.036820)+V(L_ACT1_21)*(-0.135090)+V(L_ACT1_22)*(0.056348)+V(L_ACT1_23)*(-0.176280)+V(L_ACT1_24)*(0.151111)+V(L_ACT1_25)*(0.411371)+V(L_ACT1_26)*(0.254126)+V(L_ACT1_27)*(0.272411)+V(L_ACT1_28)*(0.461332)+V(L_ACT1_29)*(0.340406)+V(L_ACT1_30)*(0.121126)+V(L_ACT1_31)*(0.326342)+V(L_ACT1_32)*(0.091787)+(0.059961))
B2_3 L2_3 0 V=(V(L_ACT1_1)*(0.421673)+V(L_ACT1_2)*(0.255010)+V(L_ACT1_3)*(-0.104441)+V(L_ACT1_4)*(0.000854)+V(L_ACT1_5)*(0.199559)+V(L_ACT1_6)*(0.278586)+V(L_ACT1_7)*(0.119897)+V(L_ACT1_8)*(0.312779)+V(L_ACT1_9)*(0.104587)+V(L_ACT1_10)*(0.226541)+V(L_ACT1_11)*(0.041246)+V(L_ACT1_12)*(0.215645)+V(L_ACT1_13)*(0.292043)+V(L_ACT1_14)*(0.029453)+V(L_ACT1_15)*(0.254115)+V(L_ACT1_16)*(0.425485)+V(L_ACT1_17)*(0.200304)+V(L_ACT1_18)*(0.222879)+V(L_ACT1_19)*(0.039393)+V(L_ACT1_20)*(-0.026011)+V(L_ACT1_21)*(-0.234794)+V(L_ACT1_22)*(0.274934)+V(L_ACT1_23)*(-0.030801)+V(L_ACT1_24)*(0.385229)+V(L_ACT1_25)*(0.254086)+V(L_ACT1_26)*(0.329515)+V(L_ACT1_27)*(-0.014621)+V(L_ACT1_28)*(0.387892)+V(L_ACT1_29)*(0.251405)+V(L_ACT1_30)*(0.281331)+V(L_ACT1_31)*(0.044941)+V(L_ACT1_32)*(0.260164)+(0.036259))
B2_4 L2_4 0 V=(V(L_ACT1_1)*(0.436904)+V(L_ACT1_2)*(0.253135)+V(L_ACT1_3)*(-0.236688)+V(L_ACT1_4)*(-0.019568)+V(L_ACT1_5)*(0.161897)+V(L_ACT1_6)*(0.291639)+V(L_ACT1_7)*(-0.100667)+V(L_ACT1_8)*(0.030223)+V(L_ACT1_9)*(0.019636)+V(L_ACT1_10)*(-0.042294)+V(L_ACT1_11)*(0.237456)+V(L_ACT1_12)*(-0.055692)+V(L_ACT1_13)*(-0.128420)+V(L_ACT1_14)*(0.157753)+V(L_ACT1_15)*(0.219080)+V(L_ACT1_16)*(0.285535)+V(L_ACT1_17)*(-0.016264)+V(L_ACT1_18)*(0.151256)+V(L_ACT1_19)*(-0.069172)+V(L_ACT1_20)*(0.255312)+V(L_ACT1_21)*(-0.206448)+V(L_ACT1_22)*(0.219978)+V(L_ACT1_23)*(0.138504)+V(L_ACT1_24)*(0.396828)+V(L_ACT1_25)*(0.067405)+V(L_ACT1_26)*(0.207178)+V(L_ACT1_27)*(0.235736)+V(L_ACT1_28)*(0.062974)+V(L_ACT1_29)*(0.284733)+V(L_ACT1_30)*(0.074773)+V(L_ACT1_31)*(0.127564)+V(L_ACT1_32)*(0.170296)+(-0.124503))
B2_5 L2_5 0 V=(V(L_ACT1_1)*(-0.519820)+V(L_ACT1_2)*(-0.078046)+V(L_ACT1_3)*(0.197488)+V(L_ACT1_4)*(0.134821)+V(L_ACT1_5)*(-0.137688)+V(L_ACT1_6)*(-0.080086)+V(L_ACT1_7)*(0.130602)+V(L_ACT1_8)*(-0.072545)+V(L_ACT1_9)*(0.003095)+V(L_ACT1_10)*(-0.181528)+V(L_ACT1_11)*(0.013982)+V(L_ACT1_12)*(-0.139001)+V(L_ACT1_13)*(0.113051)+V(L_ACT1_14)*(0.168627)+V(L_ACT1_15)*(-0.016373)+V(L_ACT1_16)*(-0.022507)+V(L_ACT1_17)*(0.087893)+V(L_ACT1_18)*(-0.136931)+V(L_ACT1_19)*(-0.042042)+V(L_ACT1_20)*(-0.065245)+V(L_ACT1_21)*(0.315252)+V(L_ACT1_22)*(-0.196943)+V(L_ACT1_23)*(0.204791)+V(L_ACT1_24)*(-0.123664)+V(L_ACT1_25)*(0.004622)+V(L_ACT1_26)*(-0.194291)+V(L_ACT1_27)*(-0.342065)+V(L_ACT1_28)*(-0.309313)+V(L_ACT1_29)*(-0.207847)+V(L_ACT1_30)*(-0.213983)+V(L_ACT1_31)*(0.106914)+V(L_ACT1_32)*(-0.024463)+(0.159825))
B2_6 L2_6 0 V=(V(L_ACT1_1)*(0.454457)+V(L_ACT1_2)*(0.143995)+V(L_ACT1_3)*(0.149878)+V(L_ACT1_4)*(-0.014341)+V(L_ACT1_5)*(0.273006)+V(L_ACT1_6)*(0.149178)+V(L_ACT1_7)*(-0.061920)+V(L_ACT1_8)*(0.054604)+V(L_ACT1_9)*(0.025957)+V(L_ACT1_10)*(0.027751)+V(L_ACT1_11)*(0.317019)+V(L_ACT1_12)*(0.316445)+V(L_ACT1_13)*(0.200801)+V(L_ACT1_14)*(0.050998)+V(L_ACT1_15)*(0.238396)+V(L_ACT1_16)*(0.180135)+V(L_ACT1_17)*(0.112504)+V(L_ACT1_18)*(0.144251)+V(L_ACT1_19)*(-0.108976)+V(L_ACT1_20)*(0.226511)+V(L_ACT1_21)*(0.001826)+V(L_ACT1_22)*(-0.038162)+V(L_ACT1_23)*(-0.225168)+V(L_ACT1_24)*(0.253185)+V(L_ACT1_25)*(0.317948)+V(L_ACT1_26)*(0.216319)+V(L_ACT1_27)*(0.263378)+V(L_ACT1_28)*(0.528740)+V(L_ACT1_29)*(0.230078)+V(L_ACT1_30)*(0.336644)+V(L_ACT1_31)*(0.279474)+V(L_ACT1_32)*(0.011594)+(0.054914))
B2_7 L2_7 0 V=(V(L_ACT1_1)*(-0.277817)+V(L_ACT1_2)*(-0.037775)+V(L_ACT1_3)*(0.207300)+V(L_ACT1_4)*(0.204926)+V(L_ACT1_5)*(-0.094955)+V(L_ACT1_6)*(-0.090642)+V(L_ACT1_7)*(0.323592)+V(L_ACT1_8)*(-0.184446)+V(L_ACT1_9)*(0.029554)+V(L_ACT1_10)*(-0.034259)+V(L_ACT1_11)*(0.086476)+V(L_ACT1_12)*(0.230525)+V(L_ACT1_13)*(-0.033043)+V(L_ACT1_14)*(0.196348)+V(L_ACT1_15)*(-0.151225)+V(L_ACT1_16)*(-0.129830)+V(L_ACT1_17)*(-0.048369)+V(L_ACT1_18)*(-0.133016)+V(L_ACT1_19)*(0.076739)+V(L_ACT1_20)*(0.008546)+V(L_ACT1_21)*(0.293961)+V(L_ACT1_22)*(-0.230297)+V(L_ACT1_23)*(0.160906)+V(L_ACT1_24)*(-0.062007)+V(L_ACT1_25)*(-0.152605)+V(L_ACT1_26)*(0.131608)+V(L_ACT1_27)*(-0.272848)+V(L_ACT1_28)*(-0.218426)+V(L_ACT1_29)*(-0.283100)+V(L_ACT1_30)*(-0.363413)+V(L_ACT1_31)*(-0.107820)+V(L_ACT1_32)*(-0.251019)+(0.029203))
B2_8 L2_8 0 V=(V(L_ACT1_1)*(-0.499393)+V(L_ACT1_2)*(-0.209863)+V(L_ACT1_3)*(0.229044)+V(L_ACT1_4)*(-0.036662)+V(L_ACT1_5)*(-0.216908)+V(L_ACT1_6)*(-0.081223)+V(L_ACT1_7)*(0.186631)+V(L_ACT1_8)*(-0.226457)+V(L_ACT1_9)*(-0.035173)+V(L_ACT1_10)*(-0.034300)+V(L_ACT1_11)*(-0.084054)+V(L_ACT1_12)*(0.174456)+V(L_ACT1_13)*(0.166640)+V(L_ACT1_14)*(-0.037028)+V(L_ACT1_15)*(-0.007816)+V(L_ACT1_16)*(-0.059755)+V(L_ACT1_17)*(0.005702)+V(L_ACT1_18)*(0.220144)+V(L_ACT1_19)*(-0.031621)+V(L_ACT1_20)*(0.152302)+V(L_ACT1_21)*(0.188611)+V(L_ACT1_22)*(0.010945)+V(L_ACT1_23)*(0.187956)+V(L_ACT1_24)*(0.110408)+V(L_ACT1_25)*(-0.040316)+V(L_ACT1_26)*(0.030480)+V(L_ACT1_27)*(-0.526112)+V(L_ACT1_28)*(-0.076988)+V(L_ACT1_29)*(-0.216628)+V(L_ACT1_30)*(-0.521296)+V(L_ACT1_31)*(0.037289)+V(L_ACT1_32)*(-0.223448)+(-0.049772))
B2_9 L2_9 0 V=(V(L_ACT1_1)*(-0.569831)+V(L_ACT1_2)*(-0.135569)+V(L_ACT1_3)*(0.208314)+V(L_ACT1_4)*(0.115522)+V(L_ACT1_5)*(-0.040774)+V(L_ACT1_6)*(-0.152223)+V(L_ACT1_7)*(0.243567)+V(L_ACT1_8)*(-0.165147)+V(L_ACT1_9)*(-0.116925)+V(L_ACT1_10)*(-0.144602)+V(L_ACT1_11)*(-0.163186)+V(L_ACT1_12)*(0.168595)+V(L_ACT1_13)*(0.003572)+V(L_ACT1_14)*(0.148279)+V(L_ACT1_15)*(-0.045484)+V(L_ACT1_16)*(-0.197602)+V(L_ACT1_17)*(-0.027718)+V(L_ACT1_18)*(0.060057)+V(L_ACT1_19)*(-0.070865)+V(L_ACT1_20)*(0.192205)+V(L_ACT1_21)*(0.111200)+V(L_ACT1_22)*(-0.176753)+V(L_ACT1_23)*(0.210591)+V(L_ACT1_24)*(-0.167227)+V(L_ACT1_25)*(-0.093995)+V(L_ACT1_26)*(-0.227974)+V(L_ACT1_27)*(-0.068557)+V(L_ACT1_28)*(-0.239977)+V(L_ACT1_29)*(-0.061432)+V(L_ACT1_30)*(-0.170131)+V(L_ACT1_31)*(0.152032)+V(L_ACT1_32)*(-0.242730)+(0.161564))
B2_10 L2_10 0 V=(V(L_ACT1_1)*(0.501889)+V(L_ACT1_2)*(0.199469)+V(L_ACT1_3)*(0.073656)+V(L_ACT1_4)*(-0.028637)+V(L_ACT1_5)*(0.131582)+V(L_ACT1_6)*(0.043960)+V(L_ACT1_7)*(0.051533)+V(L_ACT1_8)*(0.117402)+V(L_ACT1_9)*(0.315312)+V(L_ACT1_10)*(0.177621)+V(L_ACT1_11)*(0.212870)+V(L_ACT1_12)*(0.201161)+V(L_ACT1_13)*(0.185791)+V(L_ACT1_14)*(-0.109605)+V(L_ACT1_15)*(0.218067)+V(L_ACT1_16)*(0.369733)+V(L_ACT1_17)*(0.374107)+V(L_ACT1_18)*(0.408357)+V(L_ACT1_19)*(-0.238970)+V(L_ACT1_20)*(0.097190)+V(L_ACT1_21)*(0.210475)+V(L_ACT1_22)*(-0.051885)+V(L_ACT1_23)*(-0.280875)+V(L_ACT1_24)*(0.313582)+V(L_ACT1_25)*(0.118037)+V(L_ACT1_26)*(0.063043)+V(L_ACT1_27)*(0.264557)+V(L_ACT1_28)*(0.343745)+V(L_ACT1_29)*(0.383688)+V(L_ACT1_30)*(0.254880)+V(L_ACT1_31)*(0.055916)+V(L_ACT1_32)*(-0.067079)+(0.316062))
B2_11 L2_11 0 V=(V(L_ACT1_1)*(-0.574058)+V(L_ACT1_2)*(-0.244351)+V(L_ACT1_3)*(0.307773)+V(L_ACT1_4)*(0.074512)+V(L_ACT1_5)*(-0.190513)+V(L_ACT1_6)*(-0.086225)+V(L_ACT1_7)*(0.085424)+V(L_ACT1_8)*(-0.172637)+V(L_ACT1_9)*(-0.010396)+V(L_ACT1_10)*(-0.195868)+V(L_ACT1_11)*(-0.207280)+V(L_ACT1_12)*(-0.031497)+V(L_ACT1_13)*(0.009969)+V(L_ACT1_14)*(0.100006)+V(L_ACT1_15)*(-0.079631)+V(L_ACT1_16)*(0.027005)+V(L_ACT1_17)*(-0.154491)+V(L_ACT1_18)*(-0.126246)+V(L_ACT1_19)*(0.118421)+V(L_ACT1_20)*(0.183421)+V(L_ACT1_21)*(0.139781)+V(L_ACT1_22)*(-0.079454)+V(L_ACT1_23)*(0.168996)+V(L_ACT1_24)*(-0.220607)+V(L_ACT1_25)*(0.062468)+V(L_ACT1_26)*(-0.153597)+V(L_ACT1_27)*(-0.180887)+V(L_ACT1_28)*(-0.228925)+V(L_ACT1_29)*(-0.205294)+V(L_ACT1_30)*(-0.189282)+V(L_ACT1_31)*(0.158861)+V(L_ACT1_32)*(-0.174657)+(0.343677))
B2_12 L2_12 0 V=(V(L_ACT1_1)*(-0.483865)+V(L_ACT1_2)*(0.039380)+V(L_ACT1_3)*(0.221024)+V(L_ACT1_4)*(0.196059)+V(L_ACT1_5)*(-0.244206)+V(L_ACT1_6)*(-0.112923)+V(L_ACT1_7)*(0.194285)+V(L_ACT1_8)*(-0.315077)+V(L_ACT1_9)*(-0.028755)+V(L_ACT1_10)*(-0.220047)+V(L_ACT1_11)*(0.126756)+V(L_ACT1_12)*(-0.109201)+V(L_ACT1_13)*(0.024460)+V(L_ACT1_14)*(0.224156)+V(L_ACT1_15)*(-0.083991)+V(L_ACT1_16)*(-0.315993)+V(L_ACT1_17)*(-0.118516)+V(L_ACT1_18)*(-0.195170)+V(L_ACT1_19)*(-0.047701)+V(L_ACT1_20)*(0.018689)+V(L_ACT1_21)*(0.308277)+V(L_ACT1_22)*(-0.011584)+V(L_ACT1_23)*(0.289184)+V(L_ACT1_24)*(0.076121)+V(L_ACT1_25)*(-0.162575)+V(L_ACT1_26)*(-0.024138)+V(L_ACT1_27)*(-0.280006)+V(L_ACT1_28)*(-0.235452)+V(L_ACT1_29)*(-0.056170)+V(L_ACT1_30)*(-0.153845)+V(L_ACT1_31)*(0.002966)+V(L_ACT1_32)*(-0.073388)+(0.297544))
B2_13 L2_13 0 V=(V(L_ACT1_1)*(-0.350016)+V(L_ACT1_2)*(0.064434)+V(L_ACT1_3)*(0.291255)+V(L_ACT1_4)*(0.081746)+V(L_ACT1_5)*(0.019678)+V(L_ACT1_6)*(-0.088499)+V(L_ACT1_7)*(-0.068563)+V(L_ACT1_8)*(-0.065059)+V(L_ACT1_9)*(-0.149170)+V(L_ACT1_10)*(-0.208498)+V(L_ACT1_11)*(-0.153169)+V(L_ACT1_12)*(-0.023996)+V(L_ACT1_13)*(0.109946)+V(L_ACT1_14)*(-0.073502)+V(L_ACT1_15)*(0.031628)+V(L_ACT1_16)*(-0.144385)+V(L_ACT1_17)*(-0.172514)+V(L_ACT1_18)*(0.006002)+V(L_ACT1_19)*(0.254294)+V(L_ACT1_20)*(0.173919)+V(L_ACT1_21)*(0.365426)+V(L_ACT1_22)*(-0.258367)+V(L_ACT1_23)*(0.184428)+V(L_ACT1_24)*(-0.003143)+V(L_ACT1_25)*(-0.045271)+V(L_ACT1_26)*(-0.224908)+V(L_ACT1_27)*(-0.160844)+V(L_ACT1_28)*(-0.367349)+V(L_ACT1_29)*(-0.285808)+V(L_ACT1_30)*(-0.294692)+V(L_ACT1_31)*(0.000241)+V(L_ACT1_32)*(-0.301735)+(0.230787))
B2_14 L2_14 0 V=(V(L_ACT1_1)*(0.459429)+V(L_ACT1_2)*(0.253840)+V(L_ACT1_3)*(0.143025)+V(L_ACT1_4)*(-0.023055)+V(L_ACT1_5)*(0.294698)+V(L_ACT1_6)*(0.214866)+V(L_ACT1_7)*(0.039292)+V(L_ACT1_8)*(0.264265)+V(L_ACT1_9)*(0.309463)+V(L_ACT1_10)*(0.145023)+V(L_ACT1_11)*(0.344541)+V(L_ACT1_12)*(0.181320)+V(L_ACT1_13)*(0.139242)+V(L_ACT1_14)*(0.020712)+V(L_ACT1_15)*(0.149965)+V(L_ACT1_16)*(0.333541)+V(L_ACT1_17)*(0.267455)+V(L_ACT1_18)*(0.139877)+V(L_ACT1_19)*(-0.088890)+V(L_ACT1_20)*(0.239202)+V(L_ACT1_21)*(-0.083059)+V(L_ACT1_22)*(0.004500)+V(L_ACT1_23)*(-0.140665)+V(L_ACT1_24)*(0.371749)+V(L_ACT1_25)*(0.211892)+V(L_ACT1_26)*(0.147558)+V(L_ACT1_27)*(0.012668)+V(L_ACT1_28)*(0.323623)+V(L_ACT1_29)*(0.094590)+V(L_ACT1_30)*(0.274638)+V(L_ACT1_31)*(0.248097)+V(L_ACT1_32)*(0.248435)+(-0.050693))
B2_15 L2_15 0 V=(V(L_ACT1_1)*(0.525038)+V(L_ACT1_2)*(0.025944)+V(L_ACT1_3)*(0.013650)+V(L_ACT1_4)*(-0.154704)+V(L_ACT1_5)*(0.192295)+V(L_ACT1_6)*(0.211142)+V(L_ACT1_7)*(0.074959)+V(L_ACT1_8)*(0.173730)+V(L_ACT1_9)*(0.223491)+V(L_ACT1_10)*(0.089264)+V(L_ACT1_11)*(0.181082)+V(L_ACT1_12)*(0.230269)+V(L_ACT1_13)*(0.132188)+V(L_ACT1_14)*(0.148444)+V(L_ACT1_15)*(0.419765)+V(L_ACT1_16)*(0.368990)+V(L_ACT1_17)*(0.416477)+V(L_ACT1_18)*(0.389636)+V(L_ACT1_19)*(0.133680)+V(L_ACT1_20)*(0.297118)+V(L_ACT1_21)*(-0.154454)+V(L_ACT1_22)*(0.095507)+V(L_ACT1_23)*(-0.096057)+V(L_ACT1_24)*(0.391670)+V(L_ACT1_25)*(0.229832)+V(L_ACT1_26)*(0.293376)+V(L_ACT1_27)*(0.297335)+V(L_ACT1_28)*(0.280394)+V(L_ACT1_29)*(0.067254)+V(L_ACT1_30)*(0.200338)+V(L_ACT1_31)*(0.080685)+V(L_ACT1_32)*(0.260443)+(-0.039637))
B2_16 L2_16 0 V=(V(L_ACT1_1)*(0.406194)+V(L_ACT1_2)*(0.309062)+V(L_ACT1_3)*(-0.109955)+V(L_ACT1_4)*(0.188409)+V(L_ACT1_5)*(0.031761)+V(L_ACT1_6)*(0.262123)+V(L_ACT1_7)*(-0.064257)+V(L_ACT1_8)*(0.348155)+V(L_ACT1_9)*(0.102339)+V(L_ACT1_10)*(0.257701)+V(L_ACT1_11)*(-0.009261)+V(L_ACT1_12)*(0.140456)+V(L_ACT1_13)*(-0.002002)+V(L_ACT1_14)*(0.114609)+V(L_ACT1_15)*(0.224003)+V(L_ACT1_16)*(0.168431)+V(L_ACT1_17)*(0.056166)+V(L_ACT1_18)*(0.304172)+V(L_ACT1_19)*(0.017822)+V(L_ACT1_20)*(-0.085268)+V(L_ACT1_21)*(-0.246528)+V(L_ACT1_22)*(0.110594)+V(L_ACT1_23)*(-0.147009)+V(L_ACT1_24)*(0.202702)+V(L_ACT1_25)*(0.034377)+V(L_ACT1_26)*(0.005245)+V(L_ACT1_27)*(0.080447)+V(L_ACT1_28)*(0.417341)+V(L_ACT1_29)*(0.214743)+V(L_ACT1_30)*(0.295400)+V(L_ACT1_31)*(0.069929)+V(L_ACT1_32)*(0.217416)+(-0.141264))
* ACTIVATION LAYER 2: RELU
B_ACT2_1 L_ACT2_1 0 V=(IF(V(L2_1)>0,V(L2_1),0))
B_ACT2_2 L_ACT2_2 0 V=(IF(V(L2_2)>0,V(L2_2),0))
B_ACT2_3 L_ACT2_3 0 V=(IF(V(L2_3)>0,V(L2_3),0))
B_ACT2_4 L_ACT2_4 0 V=(IF(V(L2_4)>0,V(L2_4),0))
B_ACT2_5 L_ACT2_5 0 V=(IF(V(L2_5)>0,V(L2_5),0))
B_ACT2_6 L_ACT2_6 0 V=(IF(V(L2_6)>0,V(L2_6),0))
B_ACT2_7 L_ACT2_7 0 V=(IF(V(L2_7)>0,V(L2_7),0))
B_ACT2_8 L_ACT2_8 0 V=(IF(V(L2_8)>0,V(L2_8),0))
B_ACT2_9 L_ACT2_9 0 V=(IF(V(L2_9)>0,V(L2_9),0))
B_ACT2_10 L_ACT2_10 0 V=(IF(V(L2_10)>0,V(L2_10),0))
B_ACT2_11 L_ACT2_11 0 V=(IF(V(L2_11)>0,V(L2_11),0))
B_ACT2_12 L_ACT2_12 0 V=(IF(V(L2_12)>0,V(L2_12),0))
B_ACT2_13 L_ACT2_13 0 V=(IF(V(L2_13)>0,V(L2_13),0))
B_ACT2_14 L_ACT2_14 0 V=(IF(V(L2_14)>0,V(L2_14),0))
B_ACT2_15 L_ACT2_15 0 V=(IF(V(L2_15)>0,V(L2_15),0))
B_ACT2_16 L_ACT2_16 0 V=(IF(V(L2_16)>0,V(L2_16),0))
* LAYER 3: LINEAR
B3_1 L3_1 0 V=(V(L_ACT2_1)*(0.394254)+V(L_ACT2_2)*(-0.301749)+V(L_ACT2_3)*(-0.208368)+V(L_ACT2_4)*(-0.546269)+V(L_ACT2_5)*(0.248320)+V(L_ACT2_6)*(-0.326277)+V(L_ACT2_7)*(0.467181)+V(L_ACT2_8)*(0.316530)+V(L_ACT2_9)*(0.236221)+V(L_ACT2_10)*(-0.485823)+V(L_ACT2_11)*(0.378414)+V(L_ACT2_12)*(0.397559)+V(L_ACT2_13)*(0.371682)+V(L_ACT2_14)*(-0.518798)+V(L_ACT2_15)*(-0.293578)+V(L_ACT2_16)*(-0.224551)+(0.096029))
* ACTIVATION LAYER 3: SIGMOID
B_ACT3_1 L_ACT3_1 0 V=(1/(1+EXP(-V(L3_1))))
* Connect final internal node L_ACT3_1 to external output NNOUT1
B_OUT NNOUT1 0 V=V(L_ACT3_1)
.ENDS ActorSubckt